use work.graphics_pkg.all;

package enemies_pkg is    
    type enemies_rom_type is array(0 to (2**13 - 1)) of pixel_type;    
    type enemy_types is (puffpuff);
    constant MAX_ENEMIES : integer := 4;
    constant PUFFPUFF_FRAMES : enemies_rom_type := 
   (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"95",X"64",X"95",X"01",X"01",X"01",X"95",X"64",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"1b",X"1a",X"1a",X"1a",X"1b",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"bc",X"3c",X"bc",X"7d",X"bc",X"1a",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"1a",X"bc",X"1b",X"e9",X"3c",X"bc",X"1a",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"1a",X"1a",X"bc",X"bc",X"1a",X"1a",X"e9",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"01",X"1a",X"1a",X"ef",X"74",X"1a",X"1a",X"1a",X"ef",X"ef",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"1a",X"ef",X"c7",X"9a",X"93",X"1a",X"ef",X"9a",X"9a",X"ef",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"ef",X"69",X"2e",X"2e",X"2e",X"b6",X"2e",X"2e",X"2e",X"69",X"ef",X"01",X"01",
    X"01",X"01",X"01",X"ef",X"c7",X"2e",X"93",X"7d",X"ef",X"7d",X"ef",X"2e",X"9a",X"ef",X"01",X"01",
    X"01",X"01",X"9c",X"9c",X"74",X"2e",X"7d",X"7d",X"1a",X"7d",X"7d",X"2e",X"ef",X"10",X"10",X"01",
    X"01",X"01",X"9c",X"10",X"10",X"ef",X"ef",X"9c",X"2e",X"9c",X"ef",X"ef",X"d1",X"d1",X"10",X"01",
    X"01",X"01",X"01",X"9c",X"9c",X"10",X"10",X"10",X"d1",X"c9",X"c9",X"d1",X"10",X"10",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"9c",X"9c",X"10",X"2e",X"c9",X"10",X"10",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"9c",X"10",X"10",X"95",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"2e",X"95",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"64",X"95",X"95",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"1a",X"95",X"95",X"95",X"1a",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"3c",X"1b",X"1a",X"1a",X"1a",X"2e",X"1a",X"1b",X"3c",X"01",X"01",X"01",
    X"01",X"01",X"01",X"1b",X"7d",X"3c",X"1a",X"1a",X"e9",X"1a",X"1a",X"3c",X"1b",X"3c",X"01",X"01",
    X"01",X"01",X"01",X"01",X"3c",X"1b",X"7d",X"1a",X"1a",X"1a",X"1b",X"1b",X"3c",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"1b",X"3c",X"1b",X"3c",X"3c",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"95",X"64",X"95",X"01",X"01",X"01",X"95",X"64",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"95",X"01",X"1b",X"1a",X"1a",X"1a",X"95",X"1a",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"1a",X"3c",X"bc",X"bc",X"3c",X"bc",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"bc",X"1b",X"e9",X"1b",X"bc",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"1a",X"bc",X"bc",X"1a",X"1a",X"e9",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"1a",X"ef",X"74",X"1a",X"1a",X"1a",X"74",X"ef",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"ef",X"c7",X"9a",X"93",X"1a",X"ef",X"9a",X"9a",X"ef",X"1a",X"01",
    X"01",X"01",X"01",X"01",X"ef",X"69",X"2e",X"2e",X"2e",X"b6",X"2e",X"2e",X"2e",X"69",X"ef",X"01",
    X"01",X"01",X"01",X"01",X"ef",X"c7",X"2e",X"93",X"7d",X"ef",X"7d",X"ef",X"2e",X"9a",X"ef",X"01",
    X"01",X"01",X"01",X"9c",X"9c",X"74",X"2e",X"7d",X"7d",X"1a",X"7d",X"7d",X"2e",X"ef",X"10",X"10",
    X"01",X"01",X"01",X"9c",X"10",X"10",X"ef",X"ef",X"9c",X"2e",X"9c",X"ef",X"ef",X"d1",X"d1",X"10",
    X"01",X"01",X"01",X"01",X"9c",X"9c",X"10",X"10",X"10",X"d1",X"c9",X"c9",X"d1",X"10",X"10",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"9c",X"9c",X"10",X"2e",X"c9",X"10",X"10",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"9c",X"10",X"10",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"64",X"95",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"64",X"95",X"95",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"1a",X"1a",X"1b",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"3c",X"1a",X"1a",X"1a",X"2e",X"e9",X"3c",X"3c",X"1b",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1b",X"7d",X"1a",X"1a",X"e9",X"e9",X"1a",X"1b",X"1b",X"3c",X"1b",X"01",
    X"01",X"01",X"01",X"01",X"01",X"3c",X"1b",X"1a",X"1a",X"1a",X"3c",X"3c",X"3c",X"1b",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"7d",X"7d",X"1b",X"1b",X"1b",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"64",X"95",X"01",X"01",X"01",X"95",X"64",X"95",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"95",X"1a",X"1a",X"1a",X"3c",X"01",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"bc",X"1b",X"bc",X"bc",X"1b",X"1a",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"1a",X"1a",X"bc",X"3c",X"e9",X"3c",X"bc",X"1a",X"1a",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"1a",X"1a",X"1a",X"bc",X"bc",X"1a",X"1a",X"e9",X"1a",X"01",X"01",X"01",X"01",
    X"01",X"01",X"1a",X"1a",X"ef",X"74",X"1a",X"1a",X"1a",X"ef",X"ef",X"1a",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"1a",X"ef",X"c7",X"9a",X"ef",X"1a",X"ef",X"c7",X"9a",X"93",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"ef",X"69",X"2e",X"2e",X"2e",X"ef",X"2e",X"2e",X"2e",X"69",X"ef",X"01",X"01",X"01",
    X"01",X"01",X"ef",X"c7",X"2e",X"93",X"7d",X"ef",X"1b",X"74",X"2e",X"9a",X"ef",X"01",X"01",X"01",
    X"01",X"9c",X"9c",X"74",X"2e",X"7d",X"7d",X"1a",X"3c",X"7d",X"2e",X"ef",X"10",X"10",X"01",X"01",
    X"01",X"9c",X"10",X"10",X"ef",X"ef",X"9c",X"2e",X"9c",X"ef",X"ef",X"d1",X"d1",X"10",X"01",X"01",
    X"01",X"01",X"9c",X"9c",X"10",X"10",X"10",X"d1",X"c9",X"c9",X"d1",X"10",X"10",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"9c",X"9c",X"10",X"2e",X"c9",X"10",X"10",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"9c",X"10",X"10",X"64",X"95",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"64",X"2e",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"64",X"64",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"3c",X"1a",X"1a",X"95",X"95",X"95",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"3c",X"1b",X"1b",X"1a",X"1a",X"1a",X"e9",X"1a",X"1b",X"01",X"01",X"01",X"01",
    X"01",X"01",X"1b",X"7d",X"3c",X"3c",X"1a",X"1a",X"e9",X"1a",X"1a",X"3c",X"1b",X"01",X"01",X"01",
    X"01",X"01",X"01",X"3c",X"1b",X"1b",X"3c",X"1a",X"1a",X"1a",X"1b",X"3c",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"3c",X"1b",X"3c",X"1b",X"3c",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"64",X"95",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"1b",X"1a",X"95",X"2e",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"3c",X"95",X"95",X"64",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"bc",X"1b",X"bc",X"95",X"95",X"95",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"1a",X"1a",X"bc",X"bc",X"e9",X"7d",X"95",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"2e",X"74",X"1a",X"bc",X"3c",X"bc",X"1a",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"9c",X"ef",X"1b",X"69",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"9c",X"9c",X"3c",X"ef",X"9a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"9c",X"10",X"10",X"1b",X"74",X"2e",X"1a",X"1a",X"e9",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"9c",X"9c",X"c9",X"10",X"3c",X"1b",X"2e",X"ef",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"9c",X"2e",X"d1",X"d1",X"10",X"9a",X"9a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"9c",X"9c",X"10",X"d1",X"d1",X"9c",X"9c",X"1a",X"1a",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"9c",X"9c",X"9c",X"d1",X"d1",X"9c",X"1a",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"9c",X"9c",X"95",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"2e",X"95",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"3c",X"1a",X"95",X"64",X"95",X"1a",X"1b",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1b",X"7d",X"1a",X"1a",X"1a",X"2e",X"1a",X"3c",X"7d",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"3c",X"1b",X"1a",X"bc",X"1a",X"3c",X"1b",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"3c",X"1b",X"3c",X"1b",X"1b",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"64",X"95",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"1a",X"3c",X"1a",X"01",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"1b",X"1a",X"1a",X"95",X"2e",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"1a",X"bc",X"3c",X"bc",X"95",X"95",X"64",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"1a",X"1a",X"1a",X"bc",X"bc",X"e9",X"e9",X"95",X"95",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"1a",X"2e",X"74",X"1a",X"bc",X"1b",X"3c",X"1b",X"95",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"9c",X"ef",X"1b",X"69",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"9c",X"9c",X"3c",X"ef",X"9a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"9c",X"10",X"10",X"1b",X"74",X"2e",X"1a",X"1a",X"e9",X"1a",X"1a",X"1a",X"01",X"01",
    X"01",X"9c",X"9c",X"c9",X"10",X"3c",X"1b",X"2e",X"ef",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",
    X"01",X"9c",X"2e",X"d1",X"d1",X"10",X"9a",X"9a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"9c",X"9c",X"10",X"d1",X"d1",X"9c",X"9c",X"1a",X"1a",X"1a",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"9c",X"9c",X"9c",X"d1",X"d1",X"9c",X"1a",X"1a",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"9c",X"9c",X"95",X"64",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1b",X"3c",X"95",X"95",X"2e",X"64",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"3c",X"3c",X"1a",X"1a",X"95",X"95",X"95",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"1b",X"7d",X"1b",X"1a",X"e9",X"1a",X"1a",X"1a",X"3c",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"3c",X"1b",X"3c",X"1a",X"1a",X"1a",X"1b",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"3c",X"1b",X"7d",X"1b",X"3c",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"64",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"1b",X"1a",X"1a",X"95",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"1a",X"3c",X"bc",X"95",X"2e",X"95",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"bc",X"95",X"95",X"64",X"95",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"1a",X"bc",X"bc",X"95",X"95",X"95",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"2e",X"74",X"1a",X"bc",X"1b",X"95",X"1a",X"1a",X"1a",X"1a",
    X"01",X"01",X"01",X"01",X"9c",X"ef",X"1b",X"69",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",
    X"01",X"01",X"01",X"01",X"9c",X"9c",X"3c",X"ef",X"9a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",
    X"01",X"01",X"01",X"01",X"9c",X"10",X"10",X"1b",X"74",X"2e",X"1a",X"1a",X"e9",X"1a",X"1a",X"1a",
    X"01",X"01",X"01",X"9c",X"9c",X"c9",X"10",X"3c",X"1b",X"2e",X"ef",X"1a",X"1a",X"1a",X"1a",X"1a",
    X"01",X"01",X"01",X"9c",X"2e",X"d1",X"d1",X"10",X"9a",X"9a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"01",X"9c",X"9c",X"10",X"d1",X"d1",X"9c",X"9c",X"1a",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"9c",X"9c",X"9c",X"d1",X"d1",X"9c",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"95",X"9c",X"9c",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"64",X"95",X"1a",X"1b",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"1a",X"1a",X"3c",X"3c",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1b",X"1a",X"1a",X"1a",X"2e",X"1a",X"1b",X"1b",X"3c",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"3c",X"1a",X"bc",X"bc",X"3c",X"3c",X"3c",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"1b",X"3c",X"1b",X"1b",X"1b",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"95",X"64",X"95",X"01",X"01",X"01",X"95",X"64",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"1b",X"1a",X"1a",X"1a",X"3c",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"1a",X"bc",X"bc",X"bc",X"1a",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"bc",X"e9",X"e9",X"e9",X"bc",X"1a",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"1a",X"bc",X"e9",X"2e",X"e9",X"bc",X"1a",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"1a",X"1a",X"bc",X"bc",X"bc",X"1a",X"1a",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"01",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"9c",X"1a",X"1a",X"bc",X"1a",X"1a",X"1a",X"1a",X"2e",X"1a",X"1a",X"1a",X"9c",X"01",
    X"01",X"01",X"9c",X"1a",X"1a",X"bc",X"bc",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"9c",X"01",
    X"01",X"01",X"9c",X"10",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"d1",X"9c",X"01",
    X"01",X"01",X"01",X"9c",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"9c",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"1a",X"1a",X"1a",X"95",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"2e",X"95",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"64",X"95",X"95",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"3c",X"1b",X"1a",X"95",X"95",X"95",X"1a",X"1b",X"3c",X"01",X"01",X"01",
    X"01",X"01",X"01",X"1b",X"7d",X"3c",X"1a",X"1a",X"e9",X"2e",X"1a",X"3c",X"1b",X"3c",X"01",X"01",
    X"01",X"01",X"01",X"01",X"3c",X"1b",X"7d",X"1a",X"1a",X"1a",X"1b",X"1b",X"3c",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"1b",X"3c",X"1b",X"3c",X"3c",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"64",X"95",X"01",X"01",X"01",X"95",X"64",X"95",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"1b",X"01",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1b",X"1a",X"1a",X"1a",X"3c",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"bc",X"bc",X"bc",X"1a",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"bc",X"e9",X"e9",X"e9",X"bc",X"1a",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"1a",X"1a",X"bc",X"e9",X"2e",X"e9",X"bc",X"1a",X"1a",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"1a",X"1a",X"1a",X"bc",X"bc",X"bc",X"1a",X"1a",X"1a",X"01",X"01",X"01",X"01",
    X"01",X"01",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",X"01",
    X"01",X"9c",X"1a",X"1a",X"bc",X"1a",X"1a",X"1a",X"1a",X"2e",X"1a",X"1a",X"1a",X"9c",X"01",X"01",
    X"01",X"9c",X"1a",X"1a",X"bc",X"bc",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"9c",X"01",X"01",
    X"01",X"9c",X"10",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"d1",X"9c",X"01",X"01",
    X"01",X"01",X"9c",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"9c",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"1a",X"95",X"95",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"2e",X"64",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"3c",X"1a",X"95",X"64",X"64",X"95",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"3c",X"1b",X"1b",X"1a",X"1a",X"95",X"95",X"95",X"1b",X"01",X"01",X"01",X"01",
    X"01",X"01",X"1b",X"7d",X"3c",X"3c",X"1a",X"1a",X"e9",X"1a",X"1a",X"3c",X"1b",X"01",X"01",X"01",
    X"01",X"01",X"01",X"3c",X"1b",X"1b",X"3c",X"1a",X"1a",X"1a",X"1b",X"3c",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"3c",X"1b",X"3c",X"1b",X"3c",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"95",X"64",X"95",X"01",X"01",X"01",X"95",X"64",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"95",X"01",X"1b",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"3c",X"1a",X"1a",X"1a",X"1b",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"1a",X"bc",X"bc",X"bc",X"1a",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"1a",X"bc",X"e9",X"e9",X"e9",X"bc",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"bc",X"e9",X"2e",X"e9",X"bc",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"1a",X"bc",X"bc",X"bc",X"1a",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"9c",X"1a",X"1a",X"bc",X"1a",X"1a",X"1a",X"1a",X"2e",X"1a",X"1a",X"1a",X"9c",
    X"01",X"01",X"01",X"9c",X"1a",X"1a",X"bc",X"bc",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"9c",
    X"01",X"01",X"01",X"9c",X"10",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"d1",X"9c",
    X"01",X"01",X"01",X"01",X"9c",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"9c",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"1a",X"1a",X"1a",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"64",X"95",X"95",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"64",X"64",X"95",X"1a",X"1b",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"3c",X"95",X"95",X"95",X"e9",X"1a",X"3c",X"3c",X"1b",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1b",X"7d",X"1a",X"1a",X"e9",X"2e",X"1a",X"1b",X"1b",X"3c",X"1b",X"01",
    X"01",X"01",X"01",X"01",X"01",X"3c",X"1b",X"1a",X"1a",X"1a",X"3c",X"3c",X"3c",X"1b",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"7d",X"7d",X"1b",X"1b",X"1b",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"64",X"95",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"1b",X"1a",X"95",X"2e",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"3c",X"95",X"95",X"64",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"bc",X"1b",X"bc",X"95",X"95",X"95",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"1a",X"1a",X"bc",X"bc",X"e9",X"7d",X"95",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"2e",X"74",X"1a",X"bc",X"3c",X"bc",X"1a",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"9c",X"ef",X"1b",X"69",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"9c",X"9c",X"3c",X"ef",X"9a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"9c",X"10",X"10",X"1b",X"74",X"2e",X"1a",X"1a",X"e9",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"9c",X"9c",X"c9",X"10",X"3c",X"1b",X"2e",X"ef",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"9c",X"2e",X"d1",X"d1",X"10",X"9a",X"9a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"9c",X"9c",X"10",X"d1",X"d1",X"9c",X"9c",X"1a",X"1a",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"9c",X"9c",X"9c",X"d1",X"d1",X"9c",X"1a",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"9c",X"9c",X"95",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"2e",X"95",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"3c",X"1a",X"95",X"64",X"95",X"1a",X"1b",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1b",X"7d",X"1a",X"1a",X"1a",X"2e",X"1a",X"3c",X"7d",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"3c",X"1b",X"1a",X"bc",X"1a",X"3c",X"1b",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"3c",X"1b",X"3c",X"1b",X"1b",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"64",X"95",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"1a",X"3c",X"1a",X"01",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"1b",X"1a",X"1a",X"95",X"2e",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"1a",X"bc",X"3c",X"bc",X"95",X"95",X"64",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"1a",X"1a",X"1a",X"bc",X"bc",X"e9",X"e9",X"95",X"95",X"95",X"01",X"01",X"01",
    X"01",X"01",X"01",X"1a",X"2e",X"74",X"1a",X"bc",X"1b",X"3c",X"1b",X"95",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"9c",X"ef",X"1b",X"69",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"9c",X"9c",X"3c",X"ef",X"9a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"9c",X"10",X"10",X"1b",X"74",X"2e",X"1a",X"1a",X"e9",X"1a",X"1a",X"1a",X"01",X"01",
    X"01",X"9c",X"9c",X"c9",X"10",X"3c",X"1b",X"2e",X"ef",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",
    X"01",X"9c",X"2e",X"d1",X"d1",X"10",X"9a",X"9a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"9c",X"9c",X"10",X"d1",X"d1",X"9c",X"9c",X"1a",X"1a",X"1a",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"9c",X"9c",X"9c",X"d1",X"d1",X"9c",X"1a",X"1a",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"9c",X"9c",X"95",X"64",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1b",X"3c",X"95",X"95",X"2e",X"64",X"95",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"3c",X"3c",X"1a",X"1a",X"95",X"95",X"95",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"1b",X"7d",X"1b",X"1a",X"e9",X"1a",X"1a",X"1a",X"3c",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"3c",X"1b",X"3c",X"1a",X"1a",X"1a",X"1b",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"3c",X"1b",X"7d",X"1b",X"3c",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"2e",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"64",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"1b",X"1a",X"1a",X"95",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"1a",X"3c",X"bc",X"95",X"2e",X"95",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"bc",X"95",X"95",X"64",X"95",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"1a",X"bc",X"bc",X"95",X"95",X"95",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1a",X"2e",X"74",X"1a",X"bc",X"1b",X"95",X"1a",X"1a",X"1a",X"1a",
    X"01",X"01",X"01",X"01",X"9c",X"ef",X"1b",X"69",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",
    X"01",X"01",X"01",X"01",X"9c",X"9c",X"3c",X"ef",X"9a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",X"1a",
    X"01",X"01",X"01",X"01",X"9c",X"10",X"10",X"1b",X"74",X"2e",X"1a",X"1a",X"e9",X"1a",X"1a",X"1a",
    X"01",X"01",X"01",X"9c",X"9c",X"c9",X"10",X"3c",X"1b",X"2e",X"ef",X"1a",X"1a",X"1a",X"1a",X"1a",
    X"01",X"01",X"01",X"9c",X"2e",X"d1",X"d1",X"10",X"9a",X"9a",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"01",X"9c",X"9c",X"10",X"d1",X"d1",X"9c",X"9c",X"1a",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"9c",X"9c",X"9c",X"d1",X"d1",X"9c",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"95",X"9c",X"9c",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"64",X"95",X"1a",X"1b",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",X"1a",X"1a",X"3c",X"3c",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"1b",X"1a",X"1a",X"1a",X"2e",X"1a",X"1b",X"1b",X"3c",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"3c",X"1a",X"bc",X"bc",X"3c",X"3c",X"3c",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"1b",X"3c",X"1b",X"1b",X"1b",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"cf",
    X"01",X"95",X"2e",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"2e",X"95",
    X"01",X"95",X"64",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"64",X"95",
    X"01",X"95",X"95",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"95",X"95",
    X"01",X"01",X"95",X"01",X"1b",X"01",X"1a",X"1a",X"1a",X"1a",X"1a",X"01",X"1b",X"01",X"95",X"01",
    X"01",X"01",X"01",X"01",X"01",X"3c",X"1a",X"bc",X"bc",X"bc",X"1a",X"7d",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"ef",X"ef",X"1a",X"1b",X"e9",X"2e",X"bc",X"7d",X"1a",X"ef",X"ef",X"01",X"01",
    X"01",X"01",X"ef",X"9a",X"2e",X"ef",X"bc",X"e9",X"e9",X"bc",X"bc",X"ef",X"9a",X"2e",X"ef",X"01",
    X"01",X"ef",X"c7",X"3c",X"7d",X"c7",X"74",X"bc",X"bc",X"bc",X"ef",X"9a",X"7d",X"7d",X"9a",X"ef",
    X"01",X"ef",X"9a",X"1b",X"3c",X"9a",X"ef",X"bc",X"bc",X"bc",X"ef",X"9a",X"7d",X"7d",X"9a",X"ef",
    X"01",X"01",X"93",X"2e",X"9a",X"9a",X"69",X"1a",X"1a",X"1a",X"69",X"9a",X"2e",X"9a",X"ef",X"01",
    X"01",X"01",X"01",X"ef",X"b6",X"69",X"ef",X"1a",X"1a",X"1a",X"ef",X"69",X"ef",X"ef",X"01",X"01",
    X"01",X"01",X"01",X"1a",X"1a",X"1a",X"1a",X"10",X"c9",X"d1",X"1a",X"1a",X"1a",X"1a",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"1a",X"10",X"10",X"2e",X"d1",X"d1",X"1a",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"1a",X"10",X"10",X"95",X"95",X"95",X"d1",X"d1",X"1a",X"01",X"01",X"01",
    X"01",X"01",X"95",X"95",X"95",X"9c",X"9c",X"95",X"95",X"95",X"9c",X"9c",X"01",X"01",X"01",X"01",
    X"01",X"95",X"95",X"95",X"95",X"95",X"9c",X"10",X"d1",X"10",X"9c",X"01",X"01",X"01",X"01",X"01",
    X"01",X"95",X"64",X"2e",X"95",X"95",X"01",X"9c",X"9c",X"9c",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"95",X"64",X"64",X"95",X"95",X"01",X"01",X"01",X"01",X"01",X"01",X"1a",X"1a",X"1a",X"01",
    X"01",X"01",X"95",X"95",X"95",X"cf",X"3c",X"1b",X"3c",X"1b",X"3c",X"1a",X"1a",X"1a",X"1a",X"1a",
    X"01",X"01",X"3c",X"1b",X"3c",X"1b",X"1b",X"3c",X"1b",X"3c",X"1b",X"1a",X"1a",X"2e",X"e9",X"1a",
    X"01",X"1b",X"1b",X"3c",X"1b",X"3c",X"3c",X"1b",X"3c",X"1b",X"3c",X"1a",X"1a",X"e9",X"1a",X"1a",
    X"01",X"3c",X"3c",X"1b",X"3c",X"1b",X"7d",X"3c",X"1b",X"3c",X"1b",X"3c",X"1a",X"1a",X"1a",X"1b",
    X"01",X"01",X"1b",X"3c",X"1b",X"cf",X"7d",X"1b",X"3c",X"1b",X"3c",X"1b",X"3c",X"1b",X"3c",X"cf",others=>X"01"
    );
end package;