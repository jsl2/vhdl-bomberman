library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.graphics_pkg.all;
use work.levels_pkg.all;

package tileset_pkg is
    subtype tile_type is integer range 0 to 127;    
    type tileset_rom_type is array(0 to (2**15 - 1)) of pixel_type;       
                                                  
    constant CASTLE_TILESET : tileset_rom_type := 
    (X"45",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"45",
    X"45",X"e5",X"e5",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"e5",X"2e",X"45",
    X"45",X"e5",X"e5",X"83",X"83",X"45",X"45",X"45",X"45",X"45",X"45",X"83",X"83",X"e5",X"2e",X"45",
    X"45",X"e5",X"e5",X"16",X"16",X"45",X"83",X"83",X"83",X"83",X"45",X"16",X"16",X"e5",X"2e",X"45",
    X"45",X"e5",X"e5",X"16",X"16",X"45",X"16",X"16",X"16",X"16",X"45",X"16",X"16",X"e5",X"2e",X"45",
    X"45",X"e5",X"e5",X"16",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"16",X"16",X"e5",X"2e",X"45",
    X"45",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"2e",X"45",
    X"45",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"45",
    X"45",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"45",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"16",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"16",
    X"16",X"83",X"83",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"83",X"16",
    X"16",X"83",X"83",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"83",X"16",
    X"16",X"83",X"83",X"93",X"93",X"93",X"00",X"00",X"00",X"00",X"93",X"93",X"93",X"83",X"83",X"16",
    X"16",X"83",X"83",X"83",X"83",X"83",X"93",X"93",X"93",X"93",X"83",X"83",X"83",X"83",X"83",X"16",
    X"93",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"93",
    X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"34",X"34",X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",
    X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",
    X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",
    X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",
    X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",
    X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"34",X"34",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",
    X"34",X"0f",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"0f",X"34",
    X"34",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"34",
    X"34",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"34",
    X"34",X"0f",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"0f",X"34",
    X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"34",X"34",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",
    X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",
    X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",
    X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",
    X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",
    X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"34",X"34",X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",
    X"0a",X"0f",X"0a",X"0a",X"0a",X"0f",X"0f",X"0f",X"0f",X"0f",X"0f",X"0a",X"0a",X"0a",X"0f",X"0a",
    X"0f",X"0f",X"0a",X"0a",X"0f",X"0f",X"0a",X"0a",X"0a",X"0a",X"0f",X"0f",X"0a",X"0a",X"0f",X"0f",
    X"0a",X"0a",X"0a",X"0f",X"0f",X"0a",X"0a",X"0f",X"0f",X"0a",X"0a",X"0f",X"0f",X"0a",X"0a",X"0a",
    X"0a",X"0a",X"0f",X"0f",X"0a",X"0a",X"0f",X"0f",X"0f",X"0f",X"0a",X"0a",X"0f",X"0f",X"0a",X"0a",
    X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",
    X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"34",X"34",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",
    X"34",X"0f",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"0f",X"34",
    X"34",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"34",
    X"34",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"34",
    X"34",X"0f",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"0f",X"34",
    X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"34",X"34",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",
    X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",
    X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",
    X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",
    X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",
    X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"34",X"34",X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"e5",X"45",X"e5",X"e5",X"5b",X"e5",
    X"93",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"2e",
    X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"2e",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",
    X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",
    X"16",X"16",X"5b",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"16",X"16",X"16",
    X"93",X"93",X"83",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"93",X"93",X"93",X"93",
    X"45",X"45",X"83",X"e5",X"16",X"00",X"00",X"00",X"00",X"00",X"16",X"e5",X"93",X"45",X"45",X"93",
    X"16",X"16",X"83",X"e5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"e5",X"93",X"16",X"45",X"93",
    X"16",X"16",X"83",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5b",X"93",X"16",X"45",X"93",
    X"93",X"93",X"83",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5b",X"93",X"93",X"93",X"93",
    X"16",X"16",X"83",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5b",X"16",X"16",X"16",X"16",
    X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"4d",X"7b",X"7b",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",
    X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"19",X"19",X"4d",X"7b",X"4d",X"7b",X"4d",X"4d",X"19",X"19",
    X"19",X"19",X"19",X"4d",X"19",X"7b",X"4d",X"4d",X"4d",X"19",X"7b",X"19",X"4d",X"4d",X"19",X"19",
    X"19",X"19",X"4d",X"7b",X"7b",X"4d",X"19",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"19",
    X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"4d",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"4d",X"7b",X"7b",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",
    X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"19",X"19",X"4d",X"7b",X"4d",X"5b",X"2e",X"45",X"2e",X"2e",
    X"19",X"19",X"19",X"4d",X"19",X"7b",X"4d",X"4d",X"4d",X"19",X"7b",X"45",X"e5",X"e5",X"5b",X"e5",
    X"19",X"19",X"4d",X"7b",X"7b",X"4d",X"45",X"45",X"4d",X"4d",X"4d",X"45",X"e5",X"e5",X"5b",X"5b",
    X"19",X"19",X"19",X"19",X"45",X"e5",X"e5",X"e5",X"45",X"19",X"19",X"45",X"45",X"45",X"45",X"45",
    X"4d",X"4d",X"4d",X"45",X"e5",X"5b",X"e5",X"e5",X"45",X"7b",X"4d",X"93",X"93",X"93",X"93",X"00",
    X"4d",X"19",X"45",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"4d",X"4d",X"83",X"83",X"83",X"93",X"00",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",
    X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"7b",X"7b",X"4d",
    X"19",X"19",X"4d",X"4d",X"7b",X"4d",X"7b",X"4d",X"19",X"19",X"4d",X"4d",X"19",X"4d",X"4d",X"4d",
    X"19",X"19",X"4d",X"4d",X"19",X"7b",X"19",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"4d",X"19",X"4d",X"7b",X"7b",X"4d",X"19",X"19",
    X"19",X"19",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"4d",X"4d",X"7b",X"4d",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",
    X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",X"4d",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",
    X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"7b",X"7b",X"4d",
    X"2e",X"2e",X"45",X"2e",X"5b",X"4d",X"7b",X"4d",X"19",X"19",X"4d",X"4d",X"19",X"4d",X"4d",X"4d",
    X"e5",X"5b",X"e5",X"e5",X"45",X"7b",X"19",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"19",X"19",X"19",
    X"5b",X"5b",X"e5",X"e5",X"45",X"4d",X"4d",X"4d",X"45",X"45",X"4d",X"7b",X"7b",X"4d",X"19",X"19",
    X"45",X"45",X"45",X"45",X"45",X"19",X"19",X"45",X"e5",X"e5",X"e5",X"45",X"19",X"19",X"19",X"19",
    X"00",X"93",X"93",X"93",X"93",X"4d",X"7b",X"45",X"e5",X"e5",X"5b",X"e5",X"45",X"4d",X"4d",X"4d",
    X"00",X"93",X"83",X"83",X"83",X"4d",X"4d",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"45",X"19",X"4d",
    X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"4d",X"7b",X"7b",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",
    X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"19",X"19",X"4d",X"7b",X"4d",X"7b",X"4d",X"4d",X"19",X"19",
    X"19",X"19",X"19",X"4d",X"19",X"7b",X"4d",X"4d",X"4d",X"19",X"7b",X"19",X"4d",X"4d",X"19",X"19",
    X"19",X"19",X"4d",X"7b",X"7b",X"4d",X"19",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"19",
    X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"4d",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"4d",X"7b",X"7b",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",
    X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"19",X"19",X"4d",X"7b",X"4d",X"7b",X"4d",X"4d",X"19",X"19",
    X"19",X"19",X"19",X"4d",X"19",X"7b",X"4d",X"4d",X"4d",X"19",X"7b",X"19",X"4d",X"4d",X"19",X"19",
    X"19",X"19",X"4d",X"7b",X"7b",X"4d",X"19",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"19",
    X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"4d",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",
    X"7b",X"7b",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"4d",
    X"4d",X"4d",X"19",X"4d",X"4d",X"19",X"19",X"4d",X"7b",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"4d",
    X"19",X"19",X"4d",X"19",X"7b",X"4d",X"4d",X"4d",X"19",X"7b",X"19",X"4d",X"4d",X"19",X"19",X"19",
    X"19",X"19",X"19",X"4d",X"7b",X"7b",X"4d",X"19",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",
    X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"19",
    X"19",X"4d",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",
    X"7b",X"7b",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"4d",
    X"4d",X"4d",X"19",X"4d",X"4d",X"19",X"19",X"4d",X"7b",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"4d",
    X"19",X"19",X"4d",X"19",X"7b",X"4d",X"4d",X"4d",X"19",X"7b",X"19",X"4d",X"4d",X"19",X"19",X"19",
    X"19",X"19",X"19",X"4d",X"7b",X"7b",X"4d",X"19",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",
    X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"19",
    X"19",X"4d",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",
    X"83",X"93",X"16",X"83",X"93",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"45",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"93",X"83",X"83",X"16",X"45",X"93",X"45",X"16",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"83",X"83",X"16",X"83",X"16",X"45",X"93",X"16",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"5b",X"16",
    X"83",X"16",X"16",X"83",X"16",X"45",X"93",X"5b",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"5b",X"16",
    X"83",X"93",X"16",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"16",X"93",X"93",X"45",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"93",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"45",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"83",X"93",X"83",X"83",X"16",X"45",X"93",X"45",X"16",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"83",X"83",X"16",X"83",X"16",X"45",X"93",X"16",X"5b",X"83",X"45",X"e5",X"5b",X"5b",X"e5",X"16",
    X"83",X"16",X"16",X"83",X"16",X"45",X"93",X"5b",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"16",X"93",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"0a",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"16",
    X"16",X"45",X"16",X"83",X"83",X"16",X"45",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"5b",
    X"16",X"16",X"83",X"93",X"93",X"83",X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"5b",
    X"16",X"83",X"93",X"2e",X"2e",X"93",X"83",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"5b",X"5b",
    X"16",X"83",X"93",X"5b",X"5b",X"93",X"83",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"5b",X"5b",
    X"16",X"16",X"83",X"93",X"93",X"83",X"16",X"e5",X"16",X"16",X"16",X"16",X"16",X"93",X"93",X"93",
    X"16",X"45",X"16",X"83",X"83",X"16",X"45",X"16",X"83",X"83",X"83",X"83",X"83",X"83",X"00",X"00",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",X"83",X"5b",X"5b",X"5b",X"83",X"83",X"93",X"00",X"00",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"83",X"45",X"16",X"16",X"16",X"83",X"83",X"93",X"00",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"83",X"83",X"83",X"83",X"16",X"45",X"16",X"16",X"93",X"93",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"93",X"83",X"83",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"93",X"93",X"83",X"16",X"16",X"83",X"83",X"83",X"83",X"16",
    X"16",X"e5",X"5b",X"e5",X"5b",X"16",X"2e",X"93",X"19",X"93",X"93",X"4d",X"19",X"19",X"7b",X"4d",
    X"16",X"e5",X"e5",X"5b",X"5b",X"16",X"7b",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"7b",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"4d",X"4d",X"7b",
    X"16",X"e5",X"5b",X"e5",X"e5",X"16",X"2e",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",
    X"16",X"16",X"16",X"16",X"00",X"00",X"16",X"83",X"16",X"83",X"16",X"83",X"16",X"83",X"45",X"45",
    X"5b",X"5b",X"16",X"83",X"83",X"00",X"93",X"93",X"83",X"93",X"16",X"93",X"45",X"83",X"16",X"e5",
    X"5b",X"5b",X"83",X"5b",X"93",X"00",X"93",X"16",X"83",X"16",X"83",X"93",X"83",X"e5",X"83",X"83",
    X"5b",X"00",X"45",X"00",X"5b",X"83",X"00",X"16",X"83",X"16",X"83",X"83",X"5b",X"00",X"e5",X"83",
    X"5b",X"00",X"45",X"00",X"00",X"00",X"83",X"00",X"83",X"16",X"83",X"00",X"83",X"00",X"5b",X"83",
    X"00",X"00",X"83",X"83",X"00",X"00",X"16",X"83",X"16",X"83",X"45",X"16",X"00",X"83",X"00",X"93",
    X"00",X"00",X"00",X"83",X"83",X"00",X"5b",X"5b",X"83",X"5b",X"5b",X"45",X"00",X"83",X"93",X"93",
    X"00",X"83",X"00",X"00",X"16",X"5b",X"83",X"16",X"93",X"16",X"83",X"5b",X"16",X"00",X"93",X"16",
    X"00",X"83",X"83",X"00",X"45",X"16",X"16",X"5b",X"16",X"5b",X"16",X"16",X"45",X"00",X"93",X"93",
    X"00",X"00",X"00",X"00",X"83",X"00",X"5b",X"e5",X"16",X"e5",X"5b",X"00",X"83",X"00",X"83",X"00",
    X"83",X"83",X"00",X"00",X"93",X"83",X"93",X"45",X"5b",X"45",X"16",X"83",X"16",X"00",X"00",X"00",
    X"00",X"83",X"00",X"93",X"16",X"93",X"83",X"e5",X"e5",X"e5",X"93",X"16",X"5b",X"16",X"00",X"16",
    X"19",X"83",X"00",X"93",X"16",X"93",X"93",X"5b",X"5b",X"5b",X"16",X"16",X"5b",X"16",X"00",X"00",
    X"19",X"00",X"83",X"83",X"93",X"16",X"93",X"5b",X"e5",X"5b",X"16",X"5b",X"16",X"83",X"00",X"00",
    X"19",X"19",X"00",X"00",X"83",X"83",X"16",X"83",X"83",X"83",X"5b",X"93",X"83",X"00",X"00",X"19",
    X"19",X"4d",X"19",X"00",X"00",X"93",X"5b",X"16",X"83",X"16",X"e5",X"16",X"00",X"00",X"19",X"4d",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"0a",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"16",X"83",X"83",X"16",X"45",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",X"83",X"93",X"93",X"83",X"16",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"2e",X"e5",X"e5",X"83",X"93",X"2e",X"2e",X"93",X"83",X"16",
    X"93",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"83",X"93",X"5b",X"5b",X"93",X"83",X"16",
    X"00",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"e5",X"16",X"83",X"93",X"93",X"83",X"16",X"16",
    X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"16",X"45",X"16",X"83",X"83",X"16",X"45",X"16",
    X"93",X"83",X"83",X"83",X"83",X"93",X"16",X"16",X"83",X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",
    X"00",X"83",X"83",X"83",X"83",X"93",X"16",X"45",X"16",X"45",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"83",X"83",X"83",X"16",X"45",X"16",X"16",X"93",X"93",X"83",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"16",X"83",X"83",X"83",X"83",X"93",X"93",X"83",X"83",X"83",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"83",X"16",X"16",X"83",X"83",X"83",X"83",X"16",X"93",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"83",X"83",X"93",X"93",X"93",X"83",X"83",X"16",X"93",X"93",X"16",X"5b",X"e5",X"5b",X"e5",X"16",
    X"19",X"4d",X"93",X"93",X"93",X"19",X"19",X"19",X"93",X"93",X"16",X"5b",X"5b",X"e5",X"e5",X"16",
    X"19",X"19",X"4d",X"4d",X"4d",X"19",X"19",X"7b",X"4d",X"4d",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"4d",X"4d",X"7b",X"7b",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"16",X"e5",X"e5",X"5b",X"e5",X"16",
    X"7b",X"2e",X"2e",X"7b",X"7b",X"2e",X"7b",X"4d",X"4d",X"7b",X"2e",X"7b",X"7b",X"4d",X"2e",X"2e",
    X"19",X"7b",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",
    X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",
    X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",
    X"7b",X"19",X"7b",X"7b",X"7b",X"7b",X"7b",X"19",X"7b",X"7b",X"7b",X"7b",X"7b",X"7b",X"7b",X"19",
    X"2e",X"7b",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"2e",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",
    X"7b",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",
    X"4d",X"4d",X"7b",X"19",X"4d",X"7b",X"7b",X"7b",X"7b",X"7b",X"7b",X"19",X"7b",X"7b",X"7b",X"7b",
    X"4d",X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"2e",X"4d",X"19",X"19",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"2e",X"19",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"4d",X"7b",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",X"7b",X"4d",X"19",
    X"19",X"4d",X"7b",X"19",X"19",X"7b",X"19",X"19",X"19",X"19",X"4d",X"7b",X"7b",X"19",X"19",X"19",
    X"19",X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"2e",X"2e",X"7b",X"7b",X"2e",X"7b",X"4d",X"4d",X"7b",X"2e",X"7b",X"7b",X"4d",X"2e",X"2e",X"7b",
    X"7b",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",X"19",
    X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",
    X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"7b",
    X"7b",X"19",X"19",X"7b",X"7b",X"7b",X"7b",X"7b",X"19",X"7b",X"7b",X"7b",X"7b",X"7b",X"7b",X"7b",
    X"7b",X"19",X"7b",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"2e",X"19",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",
    X"2e",X"7b",X"4d",X"7b",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",
    X"2e",X"7b",X"4d",X"4d",X"7b",X"7b",X"7b",X"7b",X"7b",X"7b",X"19",X"7b",X"7b",X"7b",X"7b",X"4d",
    X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"4d",X"19",X"19",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"2e",X"19",X"19",X"4d",X"7b",X"4d",X"19",X"19",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",
    X"2e",X"19",X"4d",X"7b",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",X"7b",X"4d",
    X"4d",X"19",X"4d",X"7b",X"19",X"19",X"7b",X"19",X"19",X"19",X"19",X"4d",X"7b",X"7b",X"19",X"19",
    X"4d",X"19",X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"4d",X"7b",X"7b",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",
    X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"19",X"19",X"4d",X"7b",X"4d",X"7b",X"4d",X"4d",X"19",X"19",
    X"19",X"19",X"19",X"4d",X"19",X"7b",X"4d",X"4d",X"4d",X"19",X"7b",X"19",X"4d",X"4d",X"19",X"19",
    X"19",X"19",X"4d",X"7b",X"7b",X"4d",X"19",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"19",
    X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"e5",X"e5",X"e5",X"45",X"e5",X"e5",X"e5",X"2e",X"45",X"e5",X"e5",X"45",X"e5",X"e5",X"5b",X"e5",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"2e",X"45",X"e5",X"e5",X"e5",X"45",X"e5",X"e5",X"5b",X"5b",X"e5",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"e5",X"e5",X"e5",X"e5",X"5b",X"2e",X"45",X"e5",X"e5",X"5b",X"45",X"e5",X"5b",X"5b",X"45",
    X"16",X"2e",X"45",X"e5",X"5b",X"e5",X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",
    X"16",X"e5",X"2e",X"16",X"e5",X"45",X"83",X"5b",X"45",X"45",X"45",X"16",X"45",X"45",X"45",X"45",
    X"16",X"e5",X"2e",X"16",X"e5",X"45",X"83",X"5b",X"45",X"16",X"16",X"93",X"16",X"16",X"16",X"16",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"16",X"e5",X"5b",X"e5",X"93",X"45",X"83",X"83",X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"93",
    X"16",X"e5",X"5b",X"e5",X"2e",X"2e",X"83",X"5b",X"83",X"93",X"16",X"16",X"16",X"16",X"45",X"93",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"5b",X"93",X"16",X"16",X"16",X"16",X"45",X"93",
    X"16",X"e5",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"45",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"16",X"93",X"16",X"16",X"16",X"16",
    X"45",X"45",X"45",X"45",X"45",X"83",X"83",X"5b",X"0f",X"0f",X"0f",X"0a",X"0a",X"0a",X"0f",X"0a",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"0a",X"0f",X"0f",X"0a",X"0a",X"0f",X"0f",
    X"5b",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"0a",X"0f",X"0f",X"0a",X"0a",X"0a",
    X"e5",X"5b",X"e5",X"45",X"2e",X"45",X"83",X"93",X"45",X"93",X"45",X"0a",X"0f",X"0f",X"0a",X"0a",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"93",X"93",X"45",X"16",X"0f",X"34",X"34",X"0f",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"5b",X"93",X"45",X"16",X"83",X"0f",X"34",X"34",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"0f",X"34",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"93",X"16",X"83",X"16",X"93",X"34",
    X"16",X"e5",X"16",X"2e",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"93",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"16",X"2e",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"45",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"93",X"93",X"e5",X"5b",X"e5",X"45",X"83",X"93",X"45",X"93",X"45",X"16",X"83",X"83",X"93",X"83",
    X"2e",X"2e",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"93",X"93",X"45",X"16",X"83",X"16",X"83",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"5b",X"93",X"45",X"16",X"83",X"16",X"16",X"83",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"93",X"16",X"83",X"16",X"93",X"83",
    X"45",X"45",X"45",X"45",X"45",X"83",X"83",X"5b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"19",X"19",X"19",X"19",X"4d",X"4d",X"19",
    X"5b",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"19",X"19",X"4d",X"4d",X"19",X"19",
    X"e5",X"5b",X"e5",X"45",X"2e",X"45",X"83",X"93",X"45",X"93",X"45",X"19",X"19",X"19",X"19",X"19",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"93",X"93",X"45",X"16",X"19",X"19",X"4d",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"5b",X"93",X"45",X"16",X"83",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"93",X"16",X"83",X"16",X"93",X"19",
    X"16",X"e5",X"16",X"2e",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"93",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"16",X"2e",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"45",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"93",X"93",X"e5",X"5b",X"e5",X"45",X"83",X"93",X"45",X"93",X"45",X"16",X"83",X"83",X"93",X"83",
    X"2e",X"2e",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"93",X"93",X"45",X"16",X"83",X"16",X"83",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"5b",X"93",X"45",X"16",X"83",X"16",X"16",X"83",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"93",X"16",X"83",X"16",X"93",X"83",
    X"0a",X"0f",X"0a",X"0a",X"0a",X"0f",X"0f",X"0f",X"5b",X"83",X"83",X"45",X"45",X"45",X"45",X"45",
    X"0f",X"0f",X"0a",X"0a",X"0f",X"0f",X"0a",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"0a",X"0a",X"0a",X"0f",X"0f",X"0a",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"5b",
    X"0a",X"0a",X"0f",X"0f",X"0a",X"45",X"93",X"45",X"93",X"83",X"45",X"2e",X"45",X"e5",X"5b",X"e5",
    X"0f",X"34",X"34",X"0f",X"16",X"45",X"93",X"93",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"34",X"34",X"0f",X"83",X"16",X"45",X"93",X"5b",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"34",X"0f",X"16",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"34",X"93",X"16",X"83",X"16",X"93",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"93",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"2e",X"16",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"45",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"2e",X"16",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"93",X"83",X"83",X"16",X"45",X"93",X"45",X"93",X"83",X"45",X"e5",X"5b",X"e5",X"93",X"93",
    X"83",X"83",X"16",X"83",X"16",X"45",X"93",X"93",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"2e",X"2e",
    X"83",X"16",X"16",X"83",X"16",X"45",X"93",X"5b",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"16",X"93",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"19",X"45",X"e5",X"e5",X"e5",X"5b",X"45",X"83",X"16",X"19",X"45",X"83",X"83",X"83",X"93",X"00",
    X"19",X"93",X"5b",X"e5",X"5b",X"45",X"83",X"16",X"16",X"45",X"45",X"00",X"00",X"00",X"00",X"00",
    X"19",X"83",X"83",X"45",X"45",X"83",X"16",X"93",X"83",X"45",X"83",X"00",X"93",X"93",X"93",X"93",
    X"19",X"83",X"83",X"83",X"00",X"16",X"93",X"83",X"16",X"83",X"83",X"00",X"83",X"83",X"83",X"83",
    X"19",X"93",X"93",X"83",X"00",X"93",X"83",X"16",X"93",X"83",X"83",X"00",X"83",X"83",X"83",X"83",
    X"45",X"45",X"45",X"45",X"00",X"83",X"83",X"93",X"93",X"83",X"45",X"93",X"93",X"45",X"93",X"45",
    X"45",X"e5",X"2e",X"45",X"00",X"16",X"83",X"93",X"16",X"16",X"45",X"93",X"16",X"93",X"16",X"93",
    X"45",X"e5",X"2e",X"45",X"83",X"93",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"45",X"e5",X"2e",X"45",X"83",X"00",X"45",X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"93",X"45",
    X"5b",X"5b",X"2e",X"45",X"83",X"16",X"16",X"45",X"93",X"16",X"16",X"16",X"16",X"45",X"93",X"16",
    X"5b",X"e5",X"2e",X"45",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"5b",X"e5",X"2e",X"45",X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"45",
    X"5b",X"2e",X"2e",X"45",X"16",X"93",X"16",X"16",X"16",X"16",X"45",X"93",X"16",X"16",X"16",X"16",
    X"5b",X"45",X"45",X"45",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"83",X"93",X"93",X"83",X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"93",X"45",
    X"83",X"93",X"93",X"83",X"16",X"16",X"16",X"45",X"93",X"16",X"16",X"16",X"16",X"45",X"93",X"16",
    X"83",X"83",X"83",X"83",X"93",X"45",X"45",X"83",X"83",X"45",X"5b",X"e5",X"e5",X"e5",X"45",X"45",
    X"00",X"00",X"00",X"00",X"00",X"45",X"45",X"83",X"83",X"83",X"45",X"5b",X"e5",X"e5",X"45",X"e5",
    X"93",X"93",X"93",X"93",X"00",X"83",X"83",X"00",X"83",X"83",X"83",X"45",X"45",X"83",X"83",X"e5",
    X"83",X"83",X"83",X"93",X"00",X"83",X"83",X"83",X"00",X"83",X"83",X"00",X"83",X"83",X"83",X"e5",
    X"83",X"83",X"83",X"93",X"00",X"83",X"83",X"83",X"83",X"00",X"83",X"00",X"83",X"93",X"93",X"e5",
    X"93",X"93",X"93",X"45",X"93",X"16",X"83",X"83",X"83",X"00",X"00",X"00",X"45",X"45",X"45",X"45",
    X"45",X"93",X"16",X"16",X"16",X"16",X"16",X"93",X"83",X"00",X"83",X"00",X"45",X"2e",X"e5",X"45",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"00",X"83",X"83",X"45",X"2e",X"e5",X"45",
    X"45",X"45",X"45",X"45",X"93",X"93",X"45",X"93",X"16",X"93",X"83",X"83",X"45",X"2e",X"5b",X"5b",
    X"16",X"16",X"16",X"45",X"93",X"16",X"93",X"16",X"93",X"16",X"93",X"83",X"45",X"2e",X"e5",X"5b",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",X"45",X"2e",X"e5",X"5b",
    X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"93",X"93",X"45",X"93",X"16",X"45",X"2e",X"2e",X"5b",
    X"45",X"93",X"16",X"16",X"16",X"16",X"45",X"93",X"16",X"93",X"16",X"93",X"45",X"45",X"45",X"5b",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",X"93",X"93",X"93",
    X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"93",X"16",X"93",X"45",X"83",X"93",X"93",X"93",
    X"16",X"16",X"16",X"45",X"93",X"16",X"16",X"93",X"16",X"93",X"45",X"5b",X"45",X"93",X"93",X"93",
    X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"4d",X"7b",X"7b",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",
    X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"19",X"19",X"4d",X"7b",X"4d",X"7b",X"4d",X"4d",X"19",X"19",
    X"19",X"19",X"19",X"4d",X"19",X"7b",X"4d",X"4d",X"4d",X"19",X"7b",X"19",X"4d",X"4d",X"19",X"19",
    X"19",X"19",X"4d",X"7b",X"7b",X"4d",X"19",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"19",
    X"19",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"e5",X"e5",X"e5",X"45",X"e5",X"e5",X"e5",X"2e",X"45",X"e5",X"e5",X"45",X"e5",X"e5",X"5b",X"e5",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"2e",X"45",X"e5",X"e5",X"e5",X"45",X"e5",X"e5",X"5b",X"5b",X"e5",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"4d",X"7b",X"7b",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",
    X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"19",X"19",X"4d",X"7b",X"4d",X"7b",X"4d",X"4d",X"19",X"19",
    X"19",X"19",X"19",X"4d",X"19",X"7b",X"4d",X"4d",X"4d",X"19",X"7b",X"19",X"4d",X"4d",X"19",X"19",
    X"19",X"19",X"4d",X"7b",X"7b",X"4d",X"19",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"19",
    X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"45",X"45",X"45",X"45",X"45",X"45",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",
    X"e5",X"e5",X"e5",X"45",X"e5",X"45",X"83",X"45",X"19",X"19",X"4d",X"7b",X"4d",X"4d",X"19",X"19",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"93",X"19",X"19",X"19",X"19",X"4d",X"4d",X"19",X"19",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"93",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"5b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"19",X"19",X"19",X"19",X"19",X"19",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",
    X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",
    X"e5",X"5b",X"e5",X"e5",X"45",X"e5",X"45",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",
    X"2e",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",
    X"2e",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",X"5b",
    X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",
    X"16",X"16",X"5b",X"93",X"16",X"16",X"16",X"16",X"16",X"5b",X"93",X"16",X"16",X"16",X"16",X"16",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"4d",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"4d",
    X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"4d",
    X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"4d",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"4d",
    X"16",X"16",X"16",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"93",X"16",X"16",X"16",X"16",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"2e",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"2e",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"2e",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"2e",X"7b",X"19",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"7b",X"19",X"19",X"19",X"4d",X"4d",X"19",X"19",X"19",X"4d",
    X"16",X"5b",X"5b",X"e5",X"e5",X"16",X"7b",X"4d",X"19",X"19",X"7b",X"19",X"4d",X"19",X"4d",X"4d",
    X"16",X"e5",X"5b",X"e5",X"e5",X"16",X"7b",X"4d",X"19",X"19",X"7b",X"19",X"4d",X"19",X"4d",X"2e",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"2e",X"4d",X"19",X"19",X"2e",X"19",X"4d",X"19",X"4d",X"2e",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"19",X"19",X"19",X"19",X"4d",X"19",X"4d",X"19",X"4d",X"2e",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"7b",X"4d",X"19",X"19",X"4d",X"19",X"19",X"19",X"4d",X"7b",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",
    X"16",X"e5",X"5b",X"e5",X"5b",X"16",X"19",X"19",X"19",X"19",X"19",X"7b",X"4d",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"5b",X"5b",X"16",X"7b",X"19",X"19",X"19",X"19",X"19",X"2e",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"19",
    X"16",X"45",X"16",X"83",X"83",X"16",X"45",X"16",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"4d",X"19",X"19",X"00",X"45",X"e5",X"5b",X"16",X"5b",X"e5",X"5b",X"00",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"83",X"83",X"16",X"16",X"83",X"16",X"16",X"93",X"83",X"19",X"19",X"19",
    X"19",X"19",X"19",X"7b",X"19",X"83",X"83",X"19",X"4d",X"19",X"83",X"83",X"19",X"19",X"4d",X"19",
    X"4d",X"19",X"7b",X"4d",X"19",X"00",X"00",X"4d",X"2e",X"4d",X"00",X"00",X"19",X"19",X"7b",X"19",
    X"4d",X"7b",X"4d",X"19",X"19",X"19",X"00",X"83",X"2e",X"83",X"00",X"19",X"19",X"19",X"19",X"19",
    X"19",X"7b",X"19",X"19",X"4d",X"19",X"7b",X"4d",X"2e",X"7b",X"19",X"2e",X"7b",X"19",X"19",X"7b",
    X"4d",X"19",X"19",X"19",X"4d",X"19",X"7b",X"4d",X"7b",X"7b",X"7b",X"19",X"2e",X"2e",X"19",X"7b",
    X"4d",X"19",X"4d",X"19",X"2e",X"19",X"7b",X"2e",X"4d",X"2e",X"7b",X"19",X"2e",X"19",X"19",X"7b",
    X"4d",X"19",X"4d",X"19",X"19",X"19",X"4d",X"2e",X"4d",X"4d",X"7b",X"2e",X"2e",X"4d",X"19",X"7b",
    X"7b",X"19",X"4d",X"19",X"7b",X"19",X"4d",X"7b",X"2e",X"7b",X"2e",X"19",X"19",X"4d",X"19",X"7b",
    X"7b",X"19",X"4d",X"19",X"19",X"2e",X"4d",X"19",X"19",X"7b",X"19",X"19",X"19",X"4d",X"19",X"19",
    X"7b",X"19",X"4d",X"19",X"19",X"19",X"7b",X"4d",X"19",X"19",X"2e",X"2e",X"19",X"4d",X"19",X"19",
    X"7b",X"19",X"19",X"4d",X"19",X"19",X"7b",X"2e",X"7b",X"2e",X"2e",X"19",X"19",X"19",X"2e",X"19",
    X"4d",X"7b",X"19",X"2e",X"2e",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"19",X"19",X"4d",
    X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"2e",X"4d",X"4d",X"19",X"19",X"7b",X"7b",X"19",
    X"19",X"19",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"2e",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"2e",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",X"7b",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",X"4d",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"19",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"4d",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"7b",X"16",X"e5",X"e5",X"5b",X"5b",X"16",
    X"2e",X"19",X"19",X"4d",X"4d",X"19",X"19",X"19",X"19",X"2e",X"16",X"e5",X"e5",X"5b",X"e5",X"16",
    X"2e",X"19",X"19",X"4d",X"2e",X"19",X"19",X"19",X"4d",X"2e",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"2e",X"19",X"19",X"4d",X"2e",X"19",X"19",X"4d",X"7b",X"19",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"4d",X"19",X"19",X"19",X"2e",X"19",X"19",X"19",X"7b",X"7b",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"2e",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"19",X"19",X"19",X"4d",X"19",X"19",X"19",X"4d",X"7b",X"7b",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"7b",X"19",X"19",X"4d",X"19",X"19",X"19",X"4d",X"7b",X"4d",X"16",X"5b",X"e5",X"5b",X"e5",X"16",
    X"19",X"19",X"2e",X"4d",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"16",X"5b",X"5b",X"e5",X"e5",X"16",
    X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"4d",X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"2e",X"16",X"45",X"16",X"83",X"83",X"16",X"45",X"16",
    X"7b",X"2e",X"2e",X"7b",X"7b",X"2e",X"7b",X"4d",X"4d",X"7b",X"2e",X"7b",X"7b",X"4d",X"2e",X"2e",
    X"19",X"7b",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",
    X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",
    X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",
    X"7b",X"7b",X"7b",X"7b",X"7b",X"7b",X"7b",X"19",X"7b",X"7b",X"7b",X"7b",X"7b",X"7b",X"7b",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",
    X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",
    X"7b",X"7b",X"7b",X"19",X"7b",X"7b",X"7b",X"7b",X"7b",X"7b",X"7b",X"19",X"7b",X"7b",X"7b",X"7b",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",X"7b",X"19",
    X"19",X"4d",X"4d",X"7b",X"7b",X"4d",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"2e",X"2e",X"2e",X"7b",X"7b",X"2e",X"7b",X"2e",X"2e",X"7b",X"7b",X"4d",X"4d",X"4d",X"7b",X"7b",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",
    X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",
    X"19",X"7b",X"7b",X"7b",X"7b",X"7b",X"7b",X"19",X"19",X"7b",X"7b",X"7b",X"7b",X"7b",X"7b",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",
    X"4d",X"4d",X"4d",X"7b",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"4d",X"4d",X"4d",X"4d",
    X"7b",X"7b",X"7b",X"19",X"7b",X"7b",X"7b",X"7b",X"7b",X"7b",X"7b",X"19",X"7b",X"7b",X"7b",X"7b",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",X"7b",
    X"19",X"19",X"4d",X"4d",X"7b",X"7b",X"4d",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"7b",X"4d",X"4d",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"16",X"16",X"83",X"93",X"93",X"83",X"16",X"e5",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"16",X"83",X"93",X"2e",X"2e",X"93",X"83",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"83",X"93",X"5b",X"5b",X"93",X"83",X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"16",X"83",X"93",X"93",X"83",X"16",X"e5",X"e5",X"45",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",
    X"16",X"45",X"16",X"83",X"83",X"16",X"45",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"83",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",
    X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"0a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"16",X"16",X"83",X"16",X"16",X"16",X"16",
    X"0a",X"00",X"83",X"93",X"16",X"e5",X"83",X"00",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"0a",X"93",X"83",X"93",X"16",X"45",X"83",X"93",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"0a",X"16",X"93",X"93",X"93",X"16",X"93",X"16",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"00",
    X"0f",X"83",X"16",X"45",X"5b",X"45",X"16",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",
    X"0a",X"0f",X"00",X"83",X"83",X"00",X"0f",X"0a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"83",X"83",X"83",X"83",X"83",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"16",X"45",X"93",X"45",X"16",X"16",X"16",X"16",X"83",
    X"16",X"5b",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"16",X"93",X"45",X"16",X"93",X"93",X"16",X"83",
    X"16",X"5b",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"5b",X"93",X"45",X"16",X"93",X"93",X"16",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"83",X"83",X"83",
    X"16",X"e5",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"45",X"93",X"83",X"16",X"83",X"16",X"16",X"16",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"83",X"83",X"93",X"93",X"93",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"45",X"83",X"93",X"93",X"93",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"83",X"83",X"83",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"16",X"45",X"93",X"45",X"16",X"83",X"16",X"83",X"00",
    X"16",X"e5",X"5b",X"5b",X"e5",X"45",X"83",X"5b",X"16",X"93",X"45",X"16",X"83",X"16",X"93",X"00",
    X"16",X"e5",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"00",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"00",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"83",X"16",X"83",X"16",X"93",X"00",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"16",X"e5",X"e5",X"e5",X"e5",X"45",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"16",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"16",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"00",X"16",X"45",X"93",X"16",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"16",X"93",X"16",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"e5",X"e5",X"5b",X"5b",X"45",X"83",X"5b",X"5b",X"93",X"83",X"16",X"16",X"16",X"16",X"16",
    X"16",X"e5",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"83",X"83",X"83",X"83",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"93",X"83",X"83",X"45",X"45",X"93",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"45",X"83",X"16",X"16",X"93",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"83",X"83",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"83",X"16",X"16",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"00",X"16",X"45",X"93",X"45",X"16",X"83",X"83",X"93",X"93",
    X"16",X"5b",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"16",X"93",X"45",X"16",X"83",X"16",X"83",X"83",
    X"16",X"5b",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"5b",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"45",X"93",X"93",X"93",X"83",X"16",X"93",X"83",
    X"83",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"e5",X"e5",X"e5",X"e5",X"5b",X"2e",X"45",X"e5",X"e5",X"5b",X"45",X"e5",X"5b",X"5b",X"45",
    X"16",X"2e",X"45",X"e5",X"5b",X"e5",X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"83",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",
    X"16",X"e5",X"2e",X"16",X"e5",X"45",X"83",X"5b",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"93",
    X"16",X"e5",X"2e",X"16",X"e5",X"45",X"83",X"5b",X"45",X"93",X"83",X"83",X"83",X"83",X"83",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"83",X"83",X"16",X"16",X"16",
    X"16",X"e5",X"5b",X"e5",X"93",X"93",X"83",X"83",X"45",X"93",X"45",X"45",X"83",X"93",X"93",X"93",
    X"16",X"e5",X"5b",X"e5",X"2e",X"2e",X"83",X"5b",X"83",X"93",X"45",X"16",X"83",X"83",X"83",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"5b",X"93",X"45",X"16",X"83",X"16",X"83",X"00",
    X"16",X"e5",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"16",X"00",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"83",X"16",X"83",X"16",X"93",X"00",
    X"83",X"93",X"16",X"83",X"93",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"45",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"83",X"93",X"16",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"83",X"93",X"83",X"83",X"16",X"45",X"93",X"45",X"16",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"e5",
    X"83",X"83",X"16",X"83",X"16",X"45",X"93",X"16",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"5b",X"e5",
    X"83",X"16",X"16",X"83",X"16",X"45",X"93",X"5b",X"5b",X"83",X"16",X"16",X"16",X"16",X"16",X"16",
    X"83",X"93",X"16",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"83",X"93",X"16",X"83",X"16",X"93",X"93",X"45",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",
    X"83",X"93",X"16",X"83",X"93",X"45",X"93",X"45",X"45",X"45",X"45",X"16",X"45",X"45",X"45",X"45",
    X"83",X"93",X"16",X"83",X"45",X"45",X"93",X"16",X"16",X"16",X"16",X"93",X"16",X"16",X"16",X"16",
    X"83",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"83",X"93",X"16",X"83",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",
    X"83",X"93",X"83",X"16",X"16",X"16",X"16",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",
    X"83",X"93",X"16",X"16",X"16",X"16",X"16",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",
    X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"83",X"16",X"16",X"16",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"93",X"16",X"16",X"16",
    X"83",X"93",X"45",X"5b",X"45",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"83",X"45",X"5b",X"e5",X"2e",X"5b",X"16",X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"45",
    X"83",X"45",X"5b",X"e5",X"e5",X"2e",X"5b",X"16",X"16",X"16",X"45",X"93",X"16",X"16",X"16",X"16",
    X"5b",X"83",X"45",X"5b",X"e5",X"5b",X"2e",X"5b",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"5b",X"83",X"83",X"45",X"5b",X"e5",X"e5",X"2e",X"45",X"16",X"16",X"45",X"45",X"45",X"45",X"45",
    X"5b",X"83",X"00",X"83",X"45",X"5b",X"e5",X"45",X"83",X"16",X"16",X"45",X"5b",X"2e",X"2e",X"2e",
    X"16",X"00",X"00",X"83",X"83",X"45",X"45",X"93",X"83",X"93",X"93",X"45",X"5b",X"e5",X"e5",X"e5",
    X"16",X"83",X"00",X"93",X"83",X"83",X"83",X"93",X"83",X"45",X"45",X"45",X"5b",X"e5",X"5b",X"e5",
    X"83",X"83",X"83",X"83",X"93",X"83",X"83",X"93",X"83",X"16",X"16",X"45",X"45",X"45",X"45",X"45",
    X"83",X"83",X"83",X"16",X"83",X"16",X"83",X"93",X"83",X"5b",X"5b",X"83",X"83",X"83",X"83",X"83",
    X"83",X"83",X"83",X"93",X"16",X"83",X"83",X"93",X"83",X"e5",X"5b",X"83",X"93",X"45",X"45",X"45",
    X"83",X"83",X"83",X"93",X"93",X"45",X"83",X"83",X"5b",X"5b",X"5b",X"83",X"93",X"45",X"45",X"45",
    X"00",X"83",X"00",X"83",X"93",X"16",X"83",X"5b",X"5b",X"5b",X"5b",X"83",X"93",X"93",X"93",X"93",
    X"83",X"00",X"00",X"16",X"83",X"16",X"83",X"83",X"16",X"45",X"45",X"83",X"5b",X"5b",X"5b",X"93",
    X"83",X"00",X"00",X"93",X"16",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"5b",X"45",X"45",X"93",
    X"83",X"83",X"00",X"93",X"93",X"45",X"45",X"16",X"16",X"16",X"83",X"83",X"5b",X"45",X"45",X"93",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"5b",X"2e",X"e5",X"5b",X"45",X"93",X"93",
    X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"93",X"5b",X"2e",X"e5",X"e5",X"5b",X"45",X"93",X"93",
    X"45",X"93",X"16",X"16",X"16",X"16",X"16",X"5b",X"2e",X"5b",X"e5",X"5b",X"45",X"83",X"93",X"93",
    X"93",X"93",X"93",X"93",X"93",X"93",X"45",X"2e",X"e5",X"e5",X"5b",X"45",X"83",X"16",X"93",X"93",
    X"45",X"45",X"45",X"45",X"45",X"16",X"83",X"45",X"e5",X"5b",X"45",X"83",X"83",X"93",X"83",X"e5",
    X"2e",X"2e",X"2e",X"2e",X"45",X"16",X"83",X"93",X"45",X"45",X"83",X"83",X"83",X"93",X"83",X"45",
    X"e5",X"e5",X"e5",X"2e",X"45",X"93",X"83",X"93",X"83",X"83",X"83",X"16",X"83",X"83",X"83",X"0a",
    X"e5",X"e5",X"5b",X"2e",X"45",X"16",X"83",X"93",X"83",X"16",X"16",X"93",X"83",X"83",X"45",X"0a",
    X"45",X"45",X"45",X"45",X"45",X"16",X"83",X"93",X"83",X"93",X"93",X"93",X"83",X"45",X"45",X"45",
    X"83",X"83",X"83",X"83",X"83",X"5b",X"83",X"93",X"83",X"93",X"93",X"83",X"e5",X"e5",X"e5",X"e5",
    X"45",X"5b",X"93",X"45",X"83",X"e5",X"83",X"93",X"83",X"83",X"83",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"45",X"5b",X"93",X"45",X"83",X"2e",X"45",X"93",X"83",X"45",X"45",X"e5",X"e5",X"e5",X"5b",X"e5",
    X"93",X"93",X"93",X"93",X"83",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"45",X"83",X"83",X"83",X"83",X"16",X"16",X"16",X"16",X"16",X"16",X"e5",X"e5",X"e5",X"e5",X"45",
    X"83",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"83",X"83",X"83",X"16",X"e5",X"e5",X"e5",X"e5",X"45",
    X"83",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"83",X"83",X"83",X"16",X"e5",X"e5",X"e5",X"e5",X"45",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"e5",X"45",X"e5",X"e5",X"5b",X"e5",
    X"93",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"2e",
    X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"2e",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",
    X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",
    X"16",X"16",X"5b",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"5b",X"93",X"16",X"16",X"16",X"16",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",
    X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",
    X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"16",X"16",X"16",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"93",X"16",X"16",X"16",X"16",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"19",X"19",X"19",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"19",X"19",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"19",X"19",X"4d",X"19",X"19",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"16",X"45",X"93",X"45",X"19",X"19",X"19",X"4d",X"4d",
    X"16",X"5b",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"16",X"93",X"45",X"16",X"19",X"19",X"7b",X"7b",
    X"16",X"5b",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"5b",X"93",X"45",X"16",X"19",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"19",X"19",X"19",X"4d",
    X"16",X"e5",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"45",X"93",X"93",X"16",X"83",X"19",X"4d",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"83",X"83",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"45",X"83",X"16",X"19",X"19",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"19",X"19",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"16",X"45",X"93",X"45",X"16",X"83",X"83",X"19",X"19",
    X"16",X"e5",X"5b",X"5b",X"e5",X"45",X"83",X"5b",X"16",X"93",X"45",X"16",X"83",X"16",X"83",X"19",
    X"16",X"e5",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"5b",X"93",X"45",X"16",X"83",X"16",X"16",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"00",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"00",
    X"45",X"e5",X"e5",X"e5",X"e5",X"16",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"16",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"16",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"16",X"93",X"45",X"16",X"00",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"16",X"93",X"16",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"16",X"16",X"16",X"16",X"16",X"83",X"93",X"5b",X"5b",X"83",X"45",X"5b",X"5b",X"e5",X"e5",X"16",
    X"83",X"83",X"83",X"83",X"83",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"e5",X"16",
    X"93",X"45",X"45",X"83",X"83",X"93",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"93",X"16",X"16",X"83",X"45",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"83",X"83",X"83",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"16",X"16",X"83",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"93",X"93",X"83",X"83",X"16",X"45",X"93",X"45",X"16",X"00",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"83",X"83",X"16",X"83",X"16",X"45",X"93",X"16",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"5b",X"16",
    X"83",X"93",X"16",X"83",X"16",X"45",X"93",X"5b",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"5b",X"16",
    X"83",X"93",X"16",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"93",X"93",X"93",X"45",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"e5",X"16",
    X"0a",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"16",
    X"16",X"45",X"16",X"83",X"83",X"16",X"45",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"5b",
    X"16",X"16",X"83",X"93",X"93",X"83",X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"5b",
    X"16",X"83",X"93",X"2e",X"2e",X"93",X"83",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"5b",X"5b",
    X"16",X"83",X"93",X"5b",X"5b",X"93",X"83",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"5b",X"5b",
    X"16",X"16",X"83",X"93",X"93",X"83",X"16",X"e5",X"16",X"16",X"16",X"16",X"16",X"93",X"93",X"93",
    X"16",X"45",X"16",X"83",X"83",X"16",X"45",X"16",X"83",X"83",X"83",X"83",X"83",X"83",X"00",X"00",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",X"83",X"5b",X"5b",X"5b",X"83",X"83",X"93",X"00",X"00",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"83",X"45",X"16",X"16",X"16",X"83",X"83",X"93",X"00",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"83",X"83",X"83",X"83",X"16",X"45",X"16",X"16",X"93",X"93",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"93",X"83",X"83",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"93",X"93",X"83",X"16",X"16",X"83",X"83",X"83",X"83",X"16",
    X"16",X"e5",X"5b",X"e5",X"5b",X"16",X"2e",X"93",X"19",X"93",X"93",X"83",X"19",X"7b",X"4d",X"19",
    X"16",X"e5",X"e5",X"5b",X"5b",X"16",X"7b",X"19",X"19",X"19",X"19",X"4d",X"4d",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"2e",X"4d",X"4d",X"4d",X"19",X"19",X"4d",X"4d",X"7b",X"19",
    X"16",X"e5",X"5b",X"e5",X"e5",X"16",X"2e",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",
    X"16",X"16",X"16",X"16",X"00",X"00",X"16",X"83",X"16",X"83",X"16",X"83",X"16",X"83",X"45",X"45",
    X"5b",X"5b",X"16",X"83",X"83",X"00",X"93",X"93",X"83",X"93",X"16",X"93",X"45",X"83",X"16",X"e5",
    X"5b",X"5b",X"83",X"5b",X"93",X"00",X"93",X"16",X"83",X"16",X"83",X"93",X"83",X"e5",X"83",X"83",
    X"5b",X"00",X"45",X"00",X"5b",X"83",X"00",X"16",X"83",X"16",X"83",X"83",X"5b",X"00",X"e5",X"83",
    X"5b",X"00",X"45",X"00",X"00",X"00",X"83",X"00",X"83",X"16",X"83",X"00",X"83",X"00",X"5b",X"83",
    X"00",X"00",X"83",X"83",X"00",X"00",X"16",X"83",X"16",X"83",X"45",X"16",X"00",X"83",X"00",X"93",
    X"00",X"00",X"00",X"83",X"83",X"00",X"5b",X"5b",X"83",X"5b",X"5b",X"45",X"00",X"83",X"93",X"93",
    X"00",X"83",X"00",X"00",X"16",X"5b",X"83",X"16",X"93",X"16",X"83",X"5b",X"16",X"00",X"93",X"16",
    X"00",X"83",X"83",X"00",X"45",X"16",X"16",X"5b",X"16",X"5b",X"16",X"16",X"45",X"00",X"93",X"93",
    X"00",X"00",X"00",X"00",X"83",X"00",X"5b",X"e5",X"16",X"e5",X"5b",X"00",X"83",X"00",X"83",X"00",
    X"83",X"83",X"00",X"00",X"93",X"83",X"93",X"45",X"5b",X"45",X"16",X"83",X"16",X"00",X"00",X"00",
    X"00",X"83",X"00",X"93",X"16",X"93",X"83",X"e5",X"e5",X"e5",X"93",X"16",X"5b",X"16",X"00",X"16",
    X"83",X"83",X"00",X"93",X"16",X"93",X"93",X"5b",X"5b",X"5b",X"16",X"16",X"5b",X"16",X"00",X"00",
    X"19",X"00",X"83",X"83",X"93",X"16",X"93",X"5b",X"e5",X"5b",X"16",X"5b",X"16",X"83",X"00",X"00",
    X"19",X"19",X"00",X"00",X"83",X"83",X"16",X"83",X"83",X"83",X"5b",X"93",X"83",X"00",X"00",X"19",
    X"19",X"4d",X"19",X"00",X"00",X"93",X"5b",X"16",X"83",X"16",X"e5",X"16",X"00",X"00",X"83",X"19",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"0a",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"16",X"83",X"83",X"16",X"45",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",X"83",X"93",X"93",X"83",X"16",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"2e",X"e5",X"e5",X"83",X"93",X"2e",X"2e",X"93",X"83",X"16",
    X"93",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"83",X"93",X"5b",X"5b",X"93",X"83",X"16",
    X"00",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"e5",X"16",X"83",X"93",X"93",X"83",X"16",X"16",
    X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"16",X"45",X"16",X"83",X"83",X"16",X"45",X"16",
    X"93",X"83",X"83",X"83",X"83",X"93",X"16",X"16",X"83",X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",
    X"00",X"83",X"83",X"83",X"83",X"93",X"16",X"45",X"16",X"45",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"83",X"83",X"83",X"16",X"45",X"16",X"16",X"93",X"93",X"83",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"16",X"83",X"83",X"83",X"83",X"93",X"93",X"83",X"83",X"83",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"83",X"16",X"16",X"83",X"83",X"83",X"83",X"16",X"93",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"83",X"83",X"93",X"93",X"93",X"83",X"83",X"16",X"93",X"93",X"16",X"5b",X"e5",X"5b",X"e5",X"16",
    X"83",X"19",X"93",X"93",X"93",X"19",X"83",X"16",X"93",X"93",X"16",X"5b",X"5b",X"e5",X"e5",X"16",
    X"4d",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"19",X"7b",X"4d",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"16",X"e5",X"e5",X"5b",X"e5",X"16",
    X"7b",X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",
    X"4d",X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"4d",X"7b",X"4d",X"7b",X"4d",X"4d",X"19",X"19",
    X"7b",X"4d",X"19",X"19",X"4d",X"7b",X"19",X"19",X"4d",X"19",X"7b",X"19",X"4d",X"4d",X"19",X"19",
    X"7b",X"19",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",X"19",
    X"2e",X"7b",X"7b",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"19",
    X"2e",X"4d",X"7b",X"19",X"19",X"7b",X"19",X"19",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"7b",X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"4d",X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"4d",X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",
    X"19",X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"4d",X"4d",X"7b",X"4d",X"7b",X"4d",X"4d",X"19",X"19",
    X"2e",X"4d",X"19",X"19",X"4d",X"7b",X"19",X"4d",X"4d",X"19",X"7b",X"19",X"4d",X"4d",X"19",X"19",
    X"2e",X"19",X"7b",X"19",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",X"19",
    X"19",X"4d",X"7b",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"19",
    X"19",X"4d",X"7b",X"19",X"19",X"7b",X"19",X"4d",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"19",X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"7b",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",
    X"19",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"4d",
    X"7b",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"4d",X"7b",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"4d",
    X"2e",X"19",X"19",X"4d",X"7b",X"19",X"19",X"4d",X"19",X"7b",X"19",X"4d",X"4d",X"19",X"19",X"4d",
    X"2e",X"19",X"19",X"4d",X"7b",X"4d",X"7b",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"7b",X"19",X"7b",X"7b",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",
    X"7b",X"19",X"4d",X"7b",X"19",X"19",X"7b",X"19",X"19",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"19",
    X"4d",X"19",X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",
    X"4d",X"7b",X"4d",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",
    X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"4d",
    X"19",X"7b",X"19",X"4d",X"7b",X"19",X"4d",X"4d",X"7b",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"4d",
    X"7b",X"19",X"19",X"4d",X"7b",X"19",X"4d",X"4d",X"19",X"7b",X"19",X"4d",X"4d",X"19",X"19",X"4d",
    X"7b",X"19",X"19",X"4d",X"7b",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"2e",X"19",X"4d",X"7b",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",
    X"2e",X"19",X"4d",X"7b",X"19",X"19",X"7b",X"19",X"4d",X"4d",X"7b",X"4d",X"4d",X"19",X"19",X"19",
    X"19",X"19",X"4d",X"7b",X"19",X"4d",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",X"19",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"e5",X"16",X"83",X"93",X"93",X"83",X"16",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"83",X"93",X"2e",X"2e",X"93",X"83",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",X"83",X"93",X"5b",X"5b",X"93",X"83",X"16",
    X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"45",X"e5",X"e5",X"16",X"83",X"93",X"93",X"83",X"16",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"16",X"83",X"83",X"16",X"45",X"16",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"83",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"83",
    X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"16",X"16",X"16",X"83",X"16",X"16",X"16",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0a",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"00",X"83",X"93",X"16",X"e5",X"83",X"00",X"0a",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"83",X"93",X"16",X"e5",X"83",X"93",X"0a",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"00",X"16",X"93",X"93",X"93",X"16",X"93",X"16",X"0a",
    X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",X"83",X"16",X"45",X"5b",X"45",X"16",X"83",X"0f",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0f",X"00",X"83",X"83",X"00",X"00",X"0f",X"0a",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"e5",X"e5",X"e5",X"e5",X"5b",X"2e",X"45",X"e5",X"e5",X"5b",X"45",X"e5",X"5b",X"5b",X"45",
    X"16",X"2e",X"45",X"e5",X"5b",X"e5",X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"83",
    X"16",X"e5",X"2e",X"16",X"e5",X"45",X"83",X"5b",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"83",
    X"16",X"e5",X"2e",X"16",X"e5",X"45",X"83",X"5b",X"45",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"83",X"16",X"83",X"16",X"16",X"16",X"16",
    X"16",X"e5",X"5b",X"e5",X"93",X"45",X"83",X"83",X"45",X"83",X"45",X"83",X"93",X"93",X"93",X"93",
    X"16",X"e5",X"5b",X"e5",X"2e",X"2e",X"83",X"5b",X"83",X"83",X"45",X"16",X"83",X"83",X"83",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"5b",X"83",X"45",X"16",X"83",X"16",X"83",X"00",
    X"16",X"e5",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"45",X"83",X"45",X"16",X"83",X"16",X"93",X"00",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"83",X"83",X"16",X"83",X"16",X"93",X"83",
    X"19",X"19",X"19",X"19",X"e7",X"19",X"19",X"19",X"19",X"2e",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"e7",X"8e",X"19",X"19",X"19",X"47",X"2e",X"85",X"19",X"19",X"4d",X"4d",X"19",
    X"4d",X"4d",X"19",X"e7",X"e7",X"19",X"19",X"19",X"2e",X"85",X"2e",X"19",X"4d",X"7b",X"7b",X"4d",
    X"4d",X"4d",X"4d",X"e7",X"8e",X"e7",X"47",X"f1",X"2e",X"85",X"5b",X"e2",X"19",X"4d",X"4d",X"19",
    X"e7",X"19",X"19",X"e7",X"e7",X"8e",X"f1",X"85",X"a3",X"2e",X"5b",X"f1",X"19",X"19",X"19",X"19",
    X"8e",X"e7",X"e7",X"e7",X"8e",X"e7",X"2e",X"e2",X"be",X"47",X"2e",X"f1",X"19",X"19",X"e2",X"19",
    X"34",X"8e",X"8e",X"e7",X"e7",X"2e",X"85",X"47",X"be",X"a3",X"85",X"f1",X"19",X"e2",X"2e",X"47",
    X"c8",X"d0",X"8e",X"8e",X"c8",X"2e",X"e2",X"be",X"a3",X"5b",X"85",X"a3",X"e2",X"2e",X"5b",X"e2",
    X"e7",X"c8",X"d0",X"8e",X"c8",X"2e",X"a3",X"c8",X"47",X"85",X"f1",X"e2",X"47",X"a3",X"f1",X"47",
    X"e7",X"e7",X"d0",X"d0",X"e7",X"85",X"f1",X"e7",X"f1",X"f1",X"a3",X"47",X"be",X"47",X"f1",X"19",
    X"19",X"e7",X"e7",X"34",X"e7",X"85",X"5b",X"e7",X"f1",X"e7",X"e2",X"be",X"a3",X"f1",X"f1",X"19",
    X"19",X"19",X"e7",X"c8",X"c8",X"e7",X"85",X"f1",X"e7",X"e2",X"c8",X"a3",X"47",X"5b",X"e2",X"19",
    X"19",X"19",X"19",X"c8",X"c8",X"c8",X"e7",X"f1",X"a3",X"e7",X"47",X"e2",X"2e",X"85",X"47",X"19",
    X"e7",X"e7",X"e7",X"e7",X"c8",X"c8",X"e7",X"f1",X"e7",X"47",X"5b",X"2e",X"2e",X"a3",X"19",X"19",
    X"19",X"e7",X"e7",X"19",X"e7",X"e7",X"e7",X"f1",X"e2",X"f1",X"e2",X"e2",X"47",X"19",X"7b",X"4d",
    X"19",X"7b",X"7b",X"4d",X"e7",X"19",X"19",X"19",X"47",X"a3",X"19",X"19",X"19",X"4d",X"4d",X"19",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"45",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"00",X"16",X"45",X"93",X"45",X"16",X"83",X"83",X"93",X"83",
    X"16",X"5b",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"16",X"93",X"45",X"16",X"83",X"16",X"83",X"83",
    X"16",X"5b",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"5b",X"93",X"45",X"16",X"83",X"16",X"16",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"45",X"93",X"93",X"16",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"e5",X"e5",X"e5",X"45",X"e5",X"e5",
    X"16",X"e5",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"5b",X"45",X"e5",X"5b",X"e5",X"e5",X"e5",
    X"16",X"5b",X"e5",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"93",X"83",X"16",X"93",X"83",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"45",X"83",X"16",X"93",X"83",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"e5",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"16",X"45",X"93",X"45",X"16",X"83",X"83",X"93",X"83",
    X"e5",X"5b",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"16",X"93",X"45",X"16",X"83",X"16",X"83",X"83",
    X"16",X"16",X"16",X"16",X"16",X"16",X"83",X"5b",X"5b",X"93",X"45",X"16",X"83",X"16",X"16",X"83",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",X"45",X"93",X"93",X"16",X"83",X"16",X"93",X"83",
    X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"93",X"45",X"93",X"83",X"16",X"93",X"83",
    X"16",X"16",X"5b",X"93",X"16",X"16",X"16",X"16",X"16",X"93",X"45",X"45",X"83",X"16",X"93",X"83",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",X"16",X"93",X"83",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"45",X"83",X"16",X"93",X"83",
    X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",X"16",X"16",X"16",X"16",X"16",X"83",X"93",X"83",
    X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"93",X"83",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",
    X"16",X"16",X"16",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"93",X"16",X"16",X"16",X"83",
    X"00",X"83",X"83",X"83",X"93",X"16",X"16",X"93",X"5b",X"5b",X"93",X"93",X"93",X"93",X"93",X"83",
    X"83",X"00",X"83",X"16",X"83",X"16",X"16",X"93",X"45",X"45",X"e5",X"e5",X"93",X"5b",X"45",X"83",
    X"83",X"00",X"83",X"93",X"83",X"93",X"93",X"93",X"45",X"45",X"5b",X"5b",X"93",X"45",X"16",X"83",
    X"83",X"83",X"00",X"93",X"83",X"45",X"45",X"93",X"93",X"93",X"5b",X"5b",X"93",X"45",X"16",X"83",
    X"00",X"83",X"00",X"83",X"83",X"16",X"16",X"5b",X"5b",X"93",X"93",X"93",X"93",X"93",X"93",X"83",
    X"83",X"00",X"00",X"16",X"83",X"16",X"16",X"45",X"45",X"93",X"e5",X"e5",X"e5",X"5b",X"45",X"83",
    X"83",X"00",X"00",X"93",X"16",X"93",X"93",X"45",X"45",X"93",X"5b",X"5b",X"5b",X"45",X"16",X"83",
    X"83",X"83",X"00",X"93",X"93",X"45",X"45",X"93",X"93",X"93",X"5b",X"5b",X"5b",X"45",X"16",X"83",
    X"00",X"83",X"83",X"83",X"93",X"16",X"16",X"93",X"5b",X"5b",X"93",X"93",X"93",X"93",X"93",X"83",
    X"83",X"00",X"83",X"16",X"83",X"16",X"16",X"93",X"45",X"45",X"e5",X"e5",X"93",X"45",X"45",X"83",
    X"83",X"00",X"83",X"93",X"83",X"93",X"93",X"93",X"45",X"45",X"5b",X"5b",X"93",X"45",X"16",X"83",
    X"83",X"83",X"00",X"93",X"83",X"45",X"45",X"93",X"93",X"93",X"5b",X"5b",X"93",X"45",X"16",X"83",
    X"00",X"83",X"00",X"83",X"83",X"16",X"16",X"5b",X"5b",X"93",X"93",X"93",X"93",X"93",X"93",X"83",
    X"83",X"00",X"00",X"16",X"83",X"16",X"16",X"45",X"45",X"93",X"e5",X"e5",X"e5",X"5b",X"45",X"83",
    X"83",X"00",X"00",X"93",X"16",X"93",X"93",X"45",X"45",X"93",X"5b",X"5b",X"5b",X"45",X"16",X"83",
    X"83",X"83",X"00",X"93",X"93",X"45",X"45",X"93",X"93",X"93",X"5b",X"5b",X"5b",X"45",X"16",X"83",
    X"16",X"e5",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"45",X"93",X"16",X"e5",X"e5",X"5b",X"e5",X"45",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"16",X"e5",X"e5",X"e5",X"e5",X"45",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"16",X"e5",X"e5",X"e5",X"e5",X"45",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"00",X"16",X"45",X"93",X"16",X"e5",X"5b",X"e5",X"e5",X"45",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"16",X"93",X"16",X"e5",X"5b",X"e5",X"e5",X"45",
    X"16",X"e5",X"e5",X"5b",X"5b",X"45",X"83",X"5b",X"5b",X"93",X"16",X"e5",X"e5",X"5b",X"5b",X"45",
    X"16",X"e5",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"45",X"93",X"16",X"e5",X"e5",X"5b",X"e5",X"45",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"16",X"e5",X"e5",X"e5",X"e5",X"45",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"16",X"e5",X"5b",X"e5",X"e5",X"45",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"16",X"e5",X"e5",X"e5",X"e5",X"45",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"16",X"e5",X"e5",X"e5",X"e5",X"45",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"00",X"16",X"45",X"93",X"16",X"e5",X"5b",X"e5",X"e5",X"45",
    X"16",X"5b",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"16",X"93",X"16",X"5b",X"e5",X"5b",X"e5",X"45",
    X"16",X"5b",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"5b",X"93",X"16",X"5b",X"5b",X"e5",X"e5",X"45",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"16",X"e5",X"e5",X"e5",X"e5",X"45",
    X"16",X"e5",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"45",X"93",X"16",X"e5",X"e5",X"5b",X"e5",X"45",
    X"5b",X"e5",X"e5",X"5b",X"e5",X"5b",X"2e",X"16",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",
    X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"2e",X"16",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",
    X"5b",X"e5",X"e5",X"5b",X"e5",X"e5",X"2e",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"5b",X"5b",X"5b",X"e5",X"e5",X"e5",X"2e",X"16",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",
    X"5b",X"e5",X"5b",X"e5",X"e5",X"e5",X"2e",X"16",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",
    X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"2e",X"16",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",
    X"5b",X"e5",X"2e",X"2e",X"2e",X"2e",X"e5",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",
    X"5b",X"e5",X"e5",X"5b",X"e5",X"5b",X"2e",X"16",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",
    X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"2e",X"16",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",
    X"5b",X"e5",X"e5",X"5b",X"e5",X"e5",X"2e",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"5b",X"5b",X"5b",X"e5",X"e5",X"e5",X"2e",X"16",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",
    X"5b",X"e5",X"5b",X"e5",X"e5",X"e5",X"2e",X"16",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",
    X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"2e",X"16",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",
    X"5b",X"e5",X"2e",X"2e",X"2e",X"2e",X"e5",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",
    X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",
    X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",
    X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",
    X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",
    X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",
    X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",
    X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",
    X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",
    X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"5b",X"5b",X"e5",X"5b",X"e5",X"e5",X"5b",
    X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"5b",X"e5",X"e5",X"5b",X"e5",X"e5",X"5b",
    X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"16",X"5b",X"e5",X"e5",X"e5",X"5b",X"5b",X"5b",
    X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"16",X"5b",X"e5",X"e5",X"e5",X"5b",X"e5",X"5b",
    X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"16",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"5b",X"2e",X"2e",X"2e",X"2e",X"e5",X"5b",
    X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"5b",X"5b",X"e5",X"5b",X"e5",X"e5",X"5b",
    X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"5b",X"e5",X"e5",X"5b",X"e5",X"e5",X"5b",
    X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"16",X"5b",X"e5",X"e5",X"e5",X"5b",X"5b",X"5b",
    X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"16",X"5b",X"e5",X"e5",X"e5",X"5b",X"e5",X"5b",
    X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"16",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"5b",X"2e",X"2e",X"2e",X"2e",X"e5",X"5b",
    X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"2e",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"7b",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"7b",X"2e",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"2e",X"7b",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"7b",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"2e",X"19",
    X"16",X"5b",X"5b",X"e5",X"e5",X"16",X"7b",X"4d",X"19",X"7b",X"19",X"4d",X"19",X"4d",X"19",X"19",
    X"16",X"e5",X"5b",X"e5",X"e5",X"16",X"2e",X"7b",X"19",X"7b",X"19",X"2e",X"19",X"4d",X"2e",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"2e",X"7b",X"19",X"2e",X"19",X"2e",X"19",X"4d",X"2e",X"19",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"19",X"19",X"19",X"4d",X"19",X"4d",X"19",X"4d",X"2e",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"7b",X"4d",X"19",X"4d",X"19",X"4d",X"19",X"4d",X"7b",X"4d",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"7b",X"19",X"7b",X"19",X"19",X"4d",X"4d",X"19",X"4d",X"4d",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"2e",X"19",X"7b",X"19",X"19",X"19",X"4d",X"19",X"19",X"7b",
    X"16",X"e5",X"5b",X"e5",X"5b",X"16",X"2e",X"19",X"7b",X"19",X"4d",X"4d",X"4d",X"19",X"19",X"7b",
    X"16",X"e5",X"e5",X"5b",X"5b",X"16",X"7b",X"19",X"19",X"7b",X"19",X"7b",X"19",X"4d",X"19",X"4d",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",X"19",X"4d",X"19",X"19",X"7b",X"19",X"4d",X"19",X"4d",
    X"16",X"45",X"16",X"83",X"83",X"16",X"45",X"16",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"4d",X"19",X"19",X"00",X"45",X"e5",X"5b",X"16",X"5b",X"e5",X"5b",X"00",X"19",X"19",X"19",
    X"4d",X"19",X"19",X"19",X"83",X"83",X"16",X"16",X"83",X"16",X"16",X"93",X"83",X"19",X"19",X"19",
    X"4d",X"7b",X"19",X"19",X"19",X"83",X"83",X"19",X"4d",X"19",X"83",X"83",X"19",X"19",X"4d",X"4d",
    X"7b",X"19",X"19",X"19",X"19",X"00",X"00",X"4d",X"4d",X"4d",X"00",X"00",X"19",X"19",X"19",X"19",
    X"7b",X"19",X"19",X"4d",X"19",X"7b",X"00",X"83",X"2e",X"4d",X"00",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"7b",X"7b",X"4d",X"2e",X"7b",X"19",X"2e",X"7b",X"7b",X"7b",X"19",
    X"19",X"19",X"19",X"2e",X"19",X"19",X"7b",X"4d",X"2e",X"2e",X"2e",X"7b",X"19",X"2e",X"2e",X"4d",
    X"19",X"4d",X"19",X"2e",X"19",X"19",X"7b",X"2e",X"2e",X"2e",X"7b",X"7b",X"19",X"2e",X"19",X"7b",
    X"19",X"4d",X"19",X"19",X"19",X"4d",X"4d",X"2e",X"4d",X"4d",X"7b",X"2e",X"2e",X"2e",X"19",X"19",
    X"19",X"4d",X"19",X"7b",X"19",X"4d",X"4d",X"7b",X"7b",X"7b",X"7b",X"7b",X"19",X"19",X"19",X"19",
    X"19",X"4d",X"19",X"19",X"2e",X"4d",X"4d",X"19",X"2e",X"7b",X"2e",X"19",X"19",X"19",X"4d",X"19",
    X"19",X"4d",X"19",X"19",X"19",X"4d",X"7b",X"4d",X"19",X"19",X"19",X"2e",X"19",X"4d",X"4d",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"7b",X"2e",X"19",X"19",X"2e",X"2e",X"2e",X"19",X"19",X"19",
    X"7b",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"19",X"2e",X"4d",
    X"19",X"4d",X"2e",X"2e",X"19",X"19",X"4d",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",
    X"19",X"7b",X"4d",X"19",X"19",X"19",X"19",X"19",X"2e",X"4d",X"19",X"19",X"19",X"19",X"7b",X"7b",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"2e",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",X"19",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"19",X"7b",X"2e",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"19",X"19",X"4d",X"19",X"19",X"4d",X"19",X"19",X"4d",X"4d",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"4d",X"19",X"19",X"4d",X"19",X"7b",X"19",X"19",X"19",X"2e",X"16",X"e5",X"e5",X"5b",X"5b",X"16",
    X"19",X"2e",X"19",X"4d",X"19",X"7b",X"19",X"19",X"19",X"2e",X"16",X"e5",X"e5",X"5b",X"e5",X"16",
    X"19",X"2e",X"19",X"4d",X"19",X"2e",X"19",X"19",X"4d",X"19",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"2e",X"19",X"19",X"4d",X"19",X"2e",X"19",X"4d",X"7b",X"19",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"7b",X"4d",X"19",X"19",X"19",X"2e",X"19",X"19",X"7b",X"7b",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"4d",X"4d",X"19",X"19",X"4d",X"4d",X"19",X"19",X"4d",X"2e",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"4d",X"7b",X"2e",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"7b",X"2e",X"16",X"5b",X"e5",X"5b",X"e5",X"16",
    X"19",X"19",X"19",X"4d",X"4d",X"19",X"19",X"4d",X"2e",X"4d",X"16",X"5b",X"5b",X"e5",X"e5",X"16",
    X"4d",X"19",X"2e",X"4d",X"19",X"4d",X"4d",X"4d",X"4d",X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",
    X"7b",X"19",X"19",X"19",X"19",X"19",X"2e",X"19",X"16",X"45",X"16",X"83",X"83",X"16",X"45",X"16",
    X"45",X"45",X"e5",X"e5",X"e5",X"5b",X"45",X"83",X"83",X"45",X"45",X"93",X"83",X"83",X"83",X"83",
    X"e5",X"45",X"e5",X"e5",X"5b",X"45",X"83",X"83",X"83",X"45",X"45",X"00",X"00",X"00",X"00",X"00",
    X"e5",X"83",X"83",X"45",X"45",X"83",X"83",X"83",X"00",X"83",X"83",X"00",X"93",X"93",X"93",X"93",
    X"e5",X"83",X"83",X"83",X"00",X"83",X"83",X"00",X"83",X"83",X"83",X"00",X"93",X"83",X"83",X"83",
    X"e5",X"93",X"93",X"83",X"00",X"83",X"00",X"83",X"83",X"83",X"83",X"00",X"93",X"83",X"83",X"83",
    X"45",X"45",X"45",X"45",X"00",X"00",X"00",X"83",X"83",X"83",X"16",X"93",X"45",X"93",X"93",X"93",
    X"45",X"e5",X"2e",X"45",X"00",X"83",X"00",X"83",X"93",X"16",X"16",X"16",X"16",X"16",X"93",X"45",
    X"45",X"e5",X"2e",X"45",X"83",X"83",X"00",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"5b",X"5b",X"2e",X"45",X"83",X"83",X"93",X"16",X"93",X"45",X"93",X"93",X"45",X"45",X"45",X"45",
    X"5b",X"e5",X"2e",X"45",X"83",X"93",X"16",X"93",X"16",X"93",X"16",X"93",X"45",X"16",X"16",X"16",
    X"5b",X"e5",X"2e",X"45",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"5b",X"2e",X"2e",X"45",X"16",X"93",X"45",X"93",X"93",X"45",X"45",X"45",X"45",X"45",X"93",X"45",
    X"5b",X"45",X"45",X"45",X"93",X"16",X"93",X"16",X"93",X"45",X"16",X"16",X"16",X"16",X"93",X"45",
    X"93",X"93",X"93",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"93",X"93",X"93",X"83",X"45",X"93",X"16",X"93",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"45",
    X"93",X"93",X"93",X"45",X"5b",X"45",X"93",X"16",X"93",X"16",X"16",X"93",X"45",X"16",X"16",X"16",
    X"00",X"93",X"83",X"83",X"83",X"45",X"19",X"16",X"83",X"45",X"5b",X"e5",X"e5",X"e5",X"45",X"19",
    X"00",X"00",X"00",X"00",X"00",X"45",X"45",X"16",X"16",X"83",X"45",X"5b",X"e5",X"5b",X"93",X"19",
    X"93",X"93",X"93",X"93",X"00",X"83",X"45",X"83",X"93",X"16",X"83",X"45",X"45",X"83",X"83",X"19",
    X"83",X"83",X"83",X"83",X"00",X"83",X"83",X"16",X"83",X"93",X"16",X"00",X"83",X"83",X"83",X"19",
    X"83",X"83",X"83",X"83",X"00",X"83",X"83",X"93",X"16",X"83",X"93",X"00",X"83",X"93",X"93",X"19",
    X"45",X"93",X"45",X"93",X"93",X"45",X"83",X"93",X"93",X"83",X"83",X"00",X"45",X"45",X"45",X"45",
    X"93",X"16",X"93",X"16",X"93",X"45",X"16",X"16",X"93",X"83",X"16",X"00",X"45",X"2e",X"e5",X"45",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",X"93",X"83",X"45",X"2e",X"e5",X"45",
    X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"00",X"83",X"45",X"2e",X"e5",X"45",
    X"16",X"93",X"45",X"16",X"16",X"16",X"16",X"93",X"45",X"16",X"16",X"83",X"45",X"2e",X"5b",X"5b",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",X"45",X"2e",X"e5",X"5b",
    X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"2e",X"e5",X"5b",
    X"16",X"16",X"16",X"16",X"93",X"45",X"16",X"16",X"16",X"16",X"93",X"16",X"45",X"2e",X"2e",X"5b",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"45",X"45",X"45",X"5b",
    X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"45",X"83",X"93",X"93",X"83",
    X"16",X"93",X"45",X"16",X"16",X"16",X"16",X"93",X"45",X"16",X"16",X"16",X"83",X"93",X"93",X"83",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"93",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"45",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"16",X"45",X"93",X"45",X"16",X"83",X"83",X"93",X"83",
    X"16",X"5b",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"16",X"93",X"45",X"16",X"83",X"16",X"83",X"83",
    X"16",X"5b",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"5b",X"93",X"45",X"16",X"83",X"16",X"16",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"45",X"93",X"93",X"16",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"93",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"45",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"16",X"45",X"93",X"45",X"16",X"83",X"83",X"93",X"83",
    X"16",X"e5",X"5b",X"5b",X"e5",X"45",X"83",X"5b",X"16",X"93",X"45",X"16",X"83",X"16",X"83",X"83",
    X"16",X"e5",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"5b",X"93",X"45",X"16",X"83",X"16",X"16",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"93",X"16",X"83",X"16",X"93",X"83",
    X"19",X"19",X"7b",X"7b",X"2f",X"19",X"19",X"19",X"2f",X"2f",X"19",X"19",X"19",X"19",X"4d",X"4d",
    X"19",X"2f",X"2f",X"19",X"2f",X"2f",X"2f",X"4d",X"2f",X"4d",X"2f",X"2f",X"2f",X"19",X"19",X"7b",
    X"2f",X"2f",X"2f",X"2f",X"2f",X"2f",X"2f",X"4d",X"2f",X"2f",X"7b",X"2e",X"2e",X"2f",X"19",X"19",
    X"19",X"19",X"19",X"2f",X"2f",X"2f",X"2f",X"4d",X"2f",X"2f",X"2f",X"2f",X"2e",X"7b",X"2f",X"19",
    X"19",X"19",X"2f",X"2f",X"2f",X"2f",X"7b",X"4d",X"2f",X"2f",X"2f",X"2f",X"2f",X"7b",X"2f",X"19",
    X"19",X"2f",X"2f",X"4d",X"2f",X"7b",X"7b",X"2f",X"4d",X"2f",X"2f",X"8e",X"2f",X"4d",X"4d",X"19",
    X"2f",X"2f",X"4d",X"4d",X"2f",X"7b",X"4d",X"2f",X"4d",X"4d",X"2f",X"2f",X"8e",X"2f",X"4d",X"19",
    X"2f",X"2f",X"4d",X"7b",X"2f",X"2e",X"2f",X"2f",X"2f",X"7b",X"4d",X"2f",X"2f",X"2f",X"4d",X"2f",
    X"2f",X"4d",X"7b",X"7b",X"2f",X"2e",X"2f",X"8e",X"2f",X"7b",X"7b",X"2f",X"2f",X"2e",X"7b",X"2f",
    X"4d",X"7b",X"7b",X"2f",X"2f",X"2e",X"7b",X"2f",X"8e",X"2f",X"7b",X"4d",X"19",X"2f",X"2e",X"2f",
    X"7b",X"2f",X"2f",X"2f",X"7b",X"2f",X"2e",X"2f",X"8e",X"2f",X"2e",X"4d",X"19",X"19",X"2f",X"19",
    X"2f",X"19",X"19",X"2f",X"2f",X"7b",X"4d",X"7b",X"2f",X"2e",X"7b",X"4d",X"19",X"19",X"19",X"19",
    X"19",X"4d",X"4d",X"2f",X"7b",X"2f",X"2f",X"4d",X"2e",X"7b",X"7b",X"2f",X"19",X"19",X"4d",X"4d",
    X"4d",X"4d",X"4d",X"2f",X"2f",X"19",X"19",X"19",X"2e",X"7b",X"2e",X"19",X"19",X"4d",X"7b",X"7b",
    X"19",X"19",X"19",X"2f",X"7b",X"19",X"19",X"19",X"2f",X"2e",X"7b",X"19",X"19",X"19",X"4d",X"4d",
    X"19",X"19",X"19",X"19",X"2f",X"19",X"19",X"19",X"19",X"2e",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"7b",X"7b",X"2f",X"19",X"19",X"19",X"2f",X"2f",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",
    X"2f",X"2f",X"19",X"2f",X"2f",X"2f",X"4d",X"2f",X"4d",X"2f",X"2f",X"2f",X"19",X"19",X"7b",X"7b",
    X"2f",X"2f",X"2f",X"2f",X"2f",X"2f",X"4d",X"2f",X"2f",X"7b",X"2e",X"2e",X"2f",X"19",X"19",X"19",
    X"19",X"19",X"19",X"2f",X"2f",X"2f",X"4d",X"4d",X"2f",X"2f",X"2f",X"2e",X"7b",X"7b",X"19",X"19",
    X"19",X"19",X"19",X"2f",X"2f",X"2f",X"2f",X"7b",X"4d",X"2f",X"2f",X"2f",X"2f",X"2f",X"7b",X"2f",
    X"19",X"19",X"2f",X"2f",X"4d",X"2f",X"7b",X"7b",X"2f",X"4d",X"2f",X"2f",X"8e",X"2f",X"4d",X"4d",
    X"19",X"2f",X"2f",X"4d",X"4d",X"2f",X"7b",X"4d",X"2f",X"4d",X"4d",X"2f",X"8e",X"2f",X"2f",X"4d",
    X"19",X"2f",X"2f",X"4d",X"7b",X"2f",X"2e",X"2f",X"2f",X"7b",X"4d",X"2f",X"2f",X"2f",X"2f",X"4d",
    X"2f",X"4d",X"7b",X"7b",X"2f",X"2e",X"2f",X"8e",X"7b",X"7b",X"2f",X"2f",X"2e",X"7b",X"2f",X"19",
    X"7b",X"7b",X"2f",X"2f",X"2e",X"7b",X"2f",X"8e",X"2f",X"7b",X"4d",X"19",X"2f",X"2e",X"2f",X"19",
    X"2f",X"2f",X"2f",X"7b",X"2f",X"2e",X"2f",X"8e",X"2f",X"2e",X"4d",X"19",X"19",X"2f",X"19",X"19",
    X"19",X"19",X"2f",X"2f",X"7b",X"4d",X"7b",X"2f",X"2e",X"7b",X"4d",X"19",X"19",X"19",X"19",X"19",
    X"19",X"4d",X"4d",X"2f",X"7b",X"7b",X"2e",X"2f",X"2e",X"7b",X"7b",X"2f",X"19",X"19",X"4d",X"4d",
    X"19",X"4d",X"4d",X"4d",X"2f",X"2f",X"19",X"2e",X"2e",X"2e",X"7b",X"2e",X"19",X"19",X"4d",X"7b",
    X"19",X"19",X"19",X"19",X"2f",X"7b",X"19",X"19",X"19",X"2f",X"2e",X"7b",X"19",X"19",X"19",X"4d",
    X"19",X"19",X"19",X"19",X"19",X"2f",X"19",X"19",X"19",X"19",X"2e",X"19",X"19",X"19",X"19",X"19",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"e5",X"e5",X"e5",
    X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"45",X"e5",X"45",X"e5",X"e5",X"45",X"e5",X"e5",X"e5",X"e5",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",
    X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"16",X"16",X"16",X"83",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"83",X"16",X"16",X"16",X"16",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"00",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"00",
    X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"19",X"83",X"83",X"83",X"93",X"16",X"16",X"93",X"5b",X"5b",X"93",X"93",X"93",X"93",X"93",X"83",
    X"4d",X"83",X"83",X"16",X"83",X"16",X"16",X"93",X"45",X"45",X"e5",X"e5",X"93",X"45",X"45",X"83",
    X"19",X"7b",X"83",X"93",X"83",X"93",X"93",X"93",X"45",X"45",X"5b",X"5b",X"93",X"45",X"16",X"83",
    X"19",X"4d",X"2e",X"93",X"83",X"45",X"45",X"93",X"93",X"93",X"5b",X"5b",X"93",X"45",X"16",X"83",
    X"19",X"19",X"7b",X"2e",X"83",X"16",X"16",X"5b",X"5b",X"93",X"93",X"93",X"93",X"93",X"93",X"83",
    X"19",X"19",X"19",X"4d",X"7b",X"16",X"16",X"45",X"45",X"93",X"e5",X"e5",X"e5",X"45",X"45",X"83",
    X"19",X"19",X"19",X"4d",X"19",X"2e",X"2e",X"45",X"45",X"7b",X"5b",X"5b",X"5b",X"45",X"16",X"83",
    X"19",X"19",X"19",X"4d",X"19",X"19",X"19",X"4d",X"4d",X"7b",X"5b",X"5b",X"5b",X"45",X"16",X"83",
    X"19",X"19",X"19",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"2e",X"2e",X"2e",X"7b",X"4d",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"7b",X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"7b",X"7b",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",
    X"19",X"19",X"19",X"19",X"4d",X"4d",X"19",X"19",X"19",X"19",X"7b",X"7b",X"7b",X"7b",X"7b",X"19",
    X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"7b",X"4d",X"4d",X"19",X"4d",X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"19",
    X"19",X"19",X"19",X"19",X"19",X"7b",X"7b",X"19",X"7b",X"7b",X"4d",X"4d",X"19",X"4d",X"4d",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",X"7b",X"19",X"7b",X"7b",X"19",
    X"19",X"83",X"83",X"83",X"93",X"16",X"16",X"93",X"5b",X"5b",X"93",X"93",X"93",X"93",X"93",X"83",
    X"7b",X"83",X"83",X"16",X"83",X"16",X"16",X"93",X"45",X"45",X"e5",X"e5",X"93",X"45",X"45",X"83",
    X"7b",X"2e",X"83",X"93",X"83",X"93",X"93",X"93",X"45",X"45",X"5b",X"5b",X"93",X"45",X"16",X"83",
    X"19",X"7b",X"2e",X"93",X"83",X"45",X"45",X"93",X"93",X"93",X"5b",X"5b",X"93",X"45",X"16",X"83",
    X"19",X"19",X"7b",X"2e",X"83",X"16",X"16",X"5b",X"5b",X"93",X"93",X"93",X"93",X"93",X"93",X"83",
    X"19",X"19",X"19",X"19",X"7b",X"16",X"16",X"45",X"45",X"93",X"e5",X"e5",X"e5",X"45",X"45",X"83",
    X"19",X"19",X"19",X"19",X"4d",X"7b",X"2e",X"45",X"45",X"7b",X"5b",X"5b",X"5b",X"45",X"16",X"83",
    X"19",X"19",X"19",X"19",X"4d",X"19",X"7b",X"2e",X"7b",X"7b",X"5b",X"5b",X"5b",X"45",X"16",X"83",
    X"19",X"19",X"7b",X"19",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",X"19",X"7b",X"7b",X"2e",X"2e",
    X"19",X"19",X"19",X"19",X"7b",X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"7b",X"7b",
    X"19",X"19",X"19",X"19",X"7b",X"7b",X"7b",X"7b",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"19",
    X"19",X"19",X"19",X"4d",X"4d",X"19",X"19",X"19",X"7b",X"7b",X"7b",X"7b",X"7b",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"7b",X"4d",X"4d",X"19",X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"4d",
    X"19",X"19",X"19",X"19",X"19",X"19",X"7b",X"7b",X"19",X"7b",X"7b",X"4d",X"4d",X"19",X"4d",X"4d",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",X"7b",X"19",X"7b",X"7b",
    X"5b",X"e5",X"e5",X"5b",X"e5",X"5b",X"2e",X"16",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",
    X"5b",X"e5",X"e5",X"5b",X"5b",X"5b",X"2e",X"16",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",
    X"5b",X"e5",X"e5",X"5b",X"e5",X"5b",X"2e",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"5b",X"e5",X"5b",X"e5",X"e5",X"e5",X"2e",X"16",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",
    X"5b",X"e5",X"5b",X"e5",X"e5",X"e5",X"2e",X"16",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",
    X"5b",X"e5",X"5b",X"5b",X"5b",X"e5",X"2e",X"16",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",
    X"5b",X"e5",X"e5",X"5b",X"5b",X"e5",X"2e",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",
    X"5b",X"e5",X"e5",X"5b",X"e5",X"5b",X"2e",X"16",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",
    X"5b",X"5b",X"e5",X"e5",X"e5",X"5b",X"2e",X"16",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",
    X"5b",X"5b",X"e5",X"e5",X"e5",X"5b",X"2e",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"5b",X"5b",X"e5",X"5b",X"5b",X"5b",X"2e",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",
    X"16",X"5b",X"2e",X"93",X"5b",X"5b",X"5b",X"ad",X"ad",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"16",X"5b",X"2e",X"93",X"16",X"16",X"5b",X"ad",X"ad",X"93",X"93",X"93",X"93",X"93",X"93",X"ad",
    X"16",X"16",X"16",X"45",X"16",X"16",X"5b",X"ad",X"ad",X"93",X"93",X"93",X"93",X"93",X"ad",X"ad",
    X"16",X"16",X"45",X"45",X"45",X"16",X"5b",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"45",X"45",
    X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",
    X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",
    X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",
    X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",
    X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",
    X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",
    X"ad",X"16",X"ad",X"ad",X"ad",X"45",X"45",X"45",X"45",X"45",X"ad",X"ad",X"ad",X"16",X"16",X"16",
    X"ad",X"ad",X"45",X"45",X"ad",X"16",X"16",X"16",X"16",X"16",X"ad",X"45",X"45",X"ad",X"ad",X"16",
    X"45",X"45",X"16",X"16",X"93",X"93",X"16",X"16",X"16",X"93",X"93",X"16",X"16",X"45",X"45",X"ad",
    X"16",X"16",X"16",X"93",X"93",X"ad",X"93",X"93",X"93",X"ad",X"93",X"93",X"16",X"16",X"16",X"45",
    X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"5b",X"5b",X"e5",X"5b",X"e5",X"e5",X"5b",
    X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"5b",X"e5",X"e5",X"5b",X"e5",X"e5",X"5b",
    X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"16",X"5b",X"e5",X"e5",X"e5",X"5b",X"5b",X"5b",
    X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"16",X"5b",X"e5",X"e5",X"e5",X"5b",X"e5",X"5b",
    X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"16",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"5b",X"2e",X"2e",X"2e",X"2e",X"e5",X"5b",
    X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"5b",X"2e",X"5b",X"e5",X"e5",X"e5",X"5b",
    X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"5b",X"2e",X"e5",X"e5",X"e5",X"e5",X"5b",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"5b",X"2e",X"e5",X"5b",X"e5",X"5b",X"5b",
    X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"5b",X"e5",X"2e",X"e5",X"2e",X"e5",X"e5",
    X"ad",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"ad",X"5b",X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",
    X"ad",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"ad",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",
    X"ad",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"45",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"ad",X"5b",X"5b",X"45",X"45",X"16",X"16",X"16",
    X"0a",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"16",
    X"16",X"45",X"16",X"83",X"83",X"16",X"45",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"5b",
    X"16",X"16",X"83",X"93",X"93",X"83",X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"5b",
    X"16",X"83",X"93",X"2e",X"2e",X"93",X"83",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"5b",X"5b",
    X"16",X"83",X"93",X"5b",X"5b",X"93",X"83",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"5b",X"5b",
    X"16",X"16",X"83",X"93",X"93",X"83",X"16",X"e5",X"16",X"16",X"16",X"16",X"16",X"93",X"93",X"93",
    X"16",X"45",X"16",X"83",X"83",X"16",X"45",X"16",X"83",X"83",X"83",X"83",X"83",X"83",X"00",X"00",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",X"83",X"5b",X"5b",X"5b",X"83",X"83",X"93",X"00",X"00",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"83",X"45",X"16",X"16",X"16",X"83",X"83",X"93",X"00",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"83",X"83",X"83",X"83",X"16",X"45",X"16",X"16",X"93",X"93",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"93",X"83",X"83",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"93",X"93",X"83",X"16",X"16",X"83",X"83",X"83",X"83",X"16",
    X"16",X"e5",X"5b",X"e5",X"5b",X"16",X"2e",X"93",X"4d",X"93",X"93",X"19",X"83",X"7b",X"4d",X"93",
    X"16",X"e5",X"e5",X"5b",X"5b",X"16",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"7b",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"4d",X"7b",X"19",
    X"16",X"e5",X"5b",X"e5",X"e5",X"16",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",
    X"16",X"16",X"16",X"16",X"00",X"00",X"16",X"83",X"16",X"83",X"16",X"83",X"16",X"83",X"45",X"45",
    X"5b",X"5b",X"16",X"83",X"83",X"00",X"93",X"93",X"83",X"93",X"16",X"93",X"45",X"83",X"16",X"e5",
    X"5b",X"5b",X"83",X"5b",X"93",X"00",X"93",X"16",X"83",X"16",X"83",X"93",X"83",X"e5",X"83",X"83",
    X"5b",X"00",X"45",X"00",X"5b",X"83",X"00",X"16",X"83",X"16",X"83",X"83",X"5b",X"00",X"e5",X"83",
    X"5b",X"00",X"45",X"00",X"00",X"00",X"83",X"00",X"83",X"16",X"83",X"00",X"83",X"00",X"5b",X"83",
    X"00",X"00",X"83",X"83",X"00",X"00",X"16",X"83",X"16",X"83",X"45",X"16",X"00",X"83",X"00",X"93",
    X"00",X"00",X"00",X"83",X"83",X"00",X"5b",X"5b",X"83",X"5b",X"5b",X"45",X"00",X"83",X"93",X"93",
    X"00",X"83",X"00",X"00",X"16",X"5b",X"83",X"16",X"93",X"16",X"83",X"5b",X"16",X"00",X"93",X"16",
    X"00",X"83",X"83",X"00",X"45",X"16",X"16",X"5b",X"16",X"5b",X"16",X"16",X"45",X"00",X"93",X"93",
    X"00",X"00",X"00",X"00",X"83",X"00",X"5b",X"e5",X"16",X"e5",X"5b",X"00",X"83",X"00",X"83",X"00",
    X"83",X"83",X"00",X"00",X"93",X"83",X"93",X"45",X"5b",X"45",X"16",X"83",X"16",X"00",X"00",X"00",
    X"00",X"83",X"00",X"93",X"16",X"93",X"83",X"e5",X"e5",X"e5",X"93",X"16",X"5b",X"16",X"00",X"16",
    X"83",X"83",X"00",X"93",X"16",X"93",X"93",X"5b",X"5b",X"5b",X"16",X"16",X"5b",X"16",X"00",X"00",
    X"19",X"00",X"83",X"83",X"93",X"16",X"93",X"5b",X"e5",X"5b",X"16",X"5b",X"16",X"83",X"00",X"00",
    X"19",X"19",X"00",X"00",X"83",X"83",X"16",X"83",X"83",X"83",X"5b",X"93",X"83",X"00",X"00",X"19",
    X"19",X"4d",X"19",X"00",X"00",X"93",X"5b",X"16",X"83",X"16",X"e5",X"16",X"00",X"00",X"19",X"4d",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"0a",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"16",X"83",X"83",X"16",X"45",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",X"83",X"93",X"93",X"83",X"16",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"2e",X"e5",X"e5",X"83",X"93",X"2e",X"2e",X"93",X"83",X"16",
    X"93",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"83",X"93",X"5b",X"5b",X"93",X"83",X"16",
    X"00",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"e5",X"16",X"83",X"93",X"93",X"83",X"16",X"16",
    X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"16",X"45",X"16",X"83",X"83",X"16",X"45",X"16",
    X"93",X"83",X"83",X"83",X"83",X"93",X"16",X"16",X"83",X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",
    X"00",X"83",X"83",X"83",X"83",X"93",X"16",X"45",X"16",X"45",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"83",X"83",X"83",X"16",X"45",X"16",X"16",X"93",X"93",X"83",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"16",X"83",X"83",X"83",X"83",X"93",X"93",X"83",X"83",X"83",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"83",X"16",X"16",X"83",X"83",X"83",X"83",X"16",X"93",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"83",X"83",X"93",X"93",X"93",X"83",X"83",X"16",X"93",X"93",X"16",X"5b",X"e5",X"5b",X"e5",X"16",
    X"19",X"83",X"19",X"93",X"93",X"19",X"83",X"19",X"93",X"19",X"16",X"5b",X"5b",X"e5",X"e5",X"16",
    X"4d",X"4d",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"19",X"7b",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"19",X"19",X"4d",X"4d",X"7b",X"7b",X"4d",X"4d",X"4d",X"4d",X"16",X"e5",X"e5",X"5b",X"e5",X"16",
    X"93",X"93",X"45",X"5b",X"e5",X"2e",X"5b",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"93",X"93",X"45",X"5b",X"e5",X"e5",X"2e",X"5b",X"93",X"45",X"45",X"45",X"45",X"45",X"93",X"45",
    X"93",X"93",X"83",X"45",X"5b",X"e5",X"5b",X"2e",X"5b",X"16",X"16",X"16",X"16",X"16",X"93",X"45",
    X"93",X"93",X"16",X"83",X"45",X"5b",X"e5",X"e5",X"2e",X"45",X"93",X"93",X"93",X"93",X"93",X"93",
    X"e5",X"83",X"93",X"83",X"83",X"45",X"5b",X"e5",X"45",X"83",X"16",X"45",X"45",X"45",X"45",X"45",
    X"45",X"83",X"93",X"83",X"83",X"83",X"45",X"45",X"93",X"83",X"16",X"45",X"2e",X"2e",X"2e",X"2e",
    X"0a",X"83",X"83",X"83",X"16",X"83",X"83",X"83",X"93",X"83",X"93",X"45",X"2e",X"e5",X"e5",X"e5",
    X"0a",X"45",X"83",X"83",X"93",X"16",X"16",X"83",X"93",X"83",X"16",X"45",X"2e",X"5b",X"e5",X"e5",
    X"45",X"45",X"45",X"83",X"93",X"93",X"93",X"83",X"93",X"83",X"16",X"45",X"45",X"45",X"45",X"45",
    X"e5",X"e5",X"e5",X"e5",X"83",X"93",X"93",X"83",X"93",X"83",X"5b",X"83",X"83",X"83",X"83",X"83",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"83",X"83",X"83",X"93",X"83",X"e5",X"83",X"45",X"93",X"5b",X"45",
    X"e5",X"5b",X"e5",X"e5",X"e5",X"45",X"45",X"83",X"93",X"45",X"2e",X"83",X"45",X"93",X"5b",X"45",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"83",X"93",X"93",X"93",X"93",
    X"45",X"e5",X"e5",X"e5",X"e5",X"16",X"16",X"16",X"16",X"16",X"16",X"83",X"83",X"83",X"83",X"45",
    X"45",X"e5",X"e5",X"e5",X"e5",X"16",X"83",X"83",X"83",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"83",
    X"45",X"e5",X"e5",X"e5",X"e5",X"16",X"83",X"83",X"83",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"83",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"45",X"5b",X"45",X"93",X"83",
    X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"45",X"16",X"5b",X"2e",X"e5",X"5b",X"45",X"83",
    X"16",X"16",X"16",X"16",X"93",X"45",X"16",X"16",X"16",X"5b",X"2e",X"e5",X"e5",X"5b",X"45",X"83",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"5b",X"2e",X"5b",X"e5",X"5b",X"45",X"83",X"5b",
    X"45",X"45",X"45",X"45",X"45",X"16",X"16",X"45",X"2e",X"e5",X"e5",X"5b",X"45",X"83",X"83",X"5b",
    X"2e",X"2e",X"2e",X"5b",X"45",X"16",X"16",X"83",X"45",X"e5",X"5b",X"45",X"83",X"00",X"83",X"5b",
    X"e5",X"e5",X"e5",X"5b",X"45",X"93",X"93",X"83",X"93",X"45",X"45",X"83",X"83",X"00",X"00",X"16",
    X"e5",X"5b",X"e5",X"5b",X"45",X"45",X"45",X"83",X"93",X"83",X"83",X"83",X"93",X"00",X"83",X"16",
    X"45",X"45",X"45",X"45",X"45",X"16",X"16",X"83",X"93",X"83",X"83",X"93",X"83",X"83",X"83",X"83",
    X"83",X"83",X"83",X"83",X"83",X"5b",X"5b",X"83",X"93",X"83",X"16",X"83",X"16",X"83",X"83",X"83",
    X"45",X"45",X"45",X"93",X"83",X"5b",X"e5",X"83",X"93",X"83",X"83",X"16",X"93",X"83",X"83",X"83",
    X"45",X"45",X"45",X"93",X"83",X"5b",X"5b",X"5b",X"83",X"83",X"45",X"93",X"93",X"83",X"83",X"83",
    X"93",X"93",X"93",X"93",X"83",X"5b",X"5b",X"5b",X"5b",X"83",X"16",X"93",X"83",X"00",X"83",X"00",
    X"93",X"5b",X"5b",X"5b",X"83",X"45",X"45",X"16",X"83",X"83",X"16",X"83",X"16",X"00",X"00",X"83",
    X"93",X"45",X"45",X"5b",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"16",X"93",X"00",X"00",X"83",
    X"93",X"45",X"45",X"5b",X"83",X"83",X"16",X"16",X"16",X"45",X"45",X"93",X"93",X"00",X"83",X"83",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"e5",X"45",X"e5",X"e5",X"5b",X"e5",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"2e",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"2e",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"5b",X"5b",X"5b",X"5b",
    X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"16",X"45",X"45",X"45",X"45",
    X"16",X"16",X"5b",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"5b",X"93",X"16",X"16",X"16",X"16",
    X"4d",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",
    X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",
    X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",
    X"4d",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"16",X"16",X"16",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"93",X"16",X"16",X"16",X"16",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"45",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"45",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"45",
    X"93",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"93",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"45",
    X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"93",X"16",X"16",X"16",X"00",X"16",X"e5",X"45",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"00",X"16",X"e5",X"45",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",X"45",X"45",X"45",X"83",X"00",X"16",X"16",X"16",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"93",X"16",X"16",X"16",X"83",X"00",X"83",X"83",X"45",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"00",X"83",X"93",X"45",
    X"16",X"16",X"16",X"83",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"83",X"00",X"83",X"93",X"45",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"00",X"83",X"93",X"45",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"00",X"83",X"93",X"45",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"00",X"93",X"93",X"93",X"83",X"00",X"83",X"93",X"45",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"00",X"83",X"83",X"83",X"83",X"00",X"83",X"83",X"45",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"45",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"16",X"16",X"16",
    X"5b",X"5b",X"5b",X"5b",X"5b",X"e5",X"45",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"16",
    X"93",X"93",X"93",X"93",X"93",X"e5",X"45",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"16",X"45",X"45",X"16",X"16",X"16",
    X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"16",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"45",X"45",X"45",X"45",X"e5",X"16",X"45",X"45",X"45",X"45",X"e5",X"16",X"45",X"16",X"16",X"16",
    X"5b",X"5b",X"5b",X"5b",X"e5",X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",X"16",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"16",X"16",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"e5",X"16",X"93",X"93",X"93",X"93",X"93",X"93",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"45",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"45",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"45",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"45",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"93",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"93",
    X"45",X"e5",X"16",X"00",X"16",X"16",X"16",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"93",
    X"45",X"e5",X"16",X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"16",X"16",X"16",X"00",X"83",X"45",X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",
    X"45",X"83",X"83",X"00",X"83",X"16",X"45",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",
    X"45",X"93",X"83",X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"45",X"93",X"83",X"00",X"83",X"16",X"16",X"16",X"16",X"16",X"16",X"83",X"16",X"16",X"16",X"16",
    X"45",X"93",X"83",X"00",X"83",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"45",X"93",X"83",X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"45",X"93",X"83",X"00",X"83",X"93",X"93",X"00",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"00",
    X"45",X"83",X"83",X"00",X"83",X"83",X"83",X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",
    X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"93",X"83",X"16",X"93",X"83",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"45",X"83",X"16",X"93",X"83",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"e5",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"16",X"45",X"93",X"45",X"16",X"83",X"83",X"93",X"83",
    X"e5",X"5b",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"16",X"93",X"45",X"16",X"83",X"16",X"83",X"83",
    X"16",X"16",X"16",X"16",X"16",X"16",X"83",X"5b",X"5b",X"93",X"45",X"16",X"83",X"16",X"16",X"83",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",X"45",X"93",X"93",X"16",X"83",X"16",X"93",X"83",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"93",X"45",X"93",X"45",X"93",X"83",X"16",X"93",X"83",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"45",X"45",X"83",X"16",X"93",X"83",
    X"16",X"16",X"16",X"83",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"83",X"16",X"93",X"83",
    X"93",X"93",X"93",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",X"83",X"93",X"83",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"16",X"16",X"83",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"00",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",
    X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"00",X"83",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0a",
    X"83",X"93",X"16",X"83",X"93",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"45",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"83",X"93",X"16",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"e5",
    X"83",X"93",X"83",X"83",X"16",X"45",X"93",X"45",X"16",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"e5",
    X"83",X"83",X"16",X"83",X"16",X"45",X"93",X"16",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"5b",X"e5",
    X"83",X"16",X"16",X"83",X"16",X"45",X"93",X"5b",X"5b",X"83",X"16",X"16",X"16",X"16",X"16",X"16",
    X"83",X"93",X"16",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"83",X"93",X"16",X"83",X"16",X"93",X"93",X"45",X"93",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"83",X"93",X"16",X"83",X"93",X"45",X"93",X"45",X"93",X"16",X"16",X"16",X"16",X"16",X"16",X"16",
    X"83",X"93",X"16",X"83",X"45",X"45",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"83",X"93",X"16",X"83",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"83",X"16",X"16",X"16",
    X"83",X"93",X"83",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",X"93",X"93",X"93",
    X"83",X"16",X"16",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"00",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"83",X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"00",X"93",X"83",X"83",X"83",X"83",X"83",X"83",
    X"0a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"16",X"16",X"45",X"45",X"45",X"5b",X"5b",X"ad",X"16",X"16",X"16",X"16",X"ad",X"ad",X"45",X"16",
    X"16",X"16",X"45",X"45",X"5b",X"5b",X"5b",X"ad",X"93",X"93",X"93",X"ad",X"45",X"45",X"ad",X"93",
    X"16",X"16",X"45",X"45",X"5b",X"5b",X"5b",X"ad",X"93",X"93",X"ad",X"45",X"16",X"93",X"45",X"00",
    X"16",X"45",X"45",X"45",X"45",X"5b",X"5b",X"83",X"ad",X"ad",X"45",X"16",X"16",X"93",X"00",X"00",
    X"16",X"16",X"16",X"45",X"45",X"5b",X"5b",X"83",X"16",X"ad",X"45",X"16",X"93",X"00",X"00",X"00",
    X"16",X"16",X"45",X"45",X"45",X"45",X"5b",X"83",X"ad",X"45",X"16",X"16",X"93",X"00",X"00",X"00",
    X"16",X"16",X"16",X"16",X"16",X"45",X"45",X"83",X"ad",X"45",X"16",X"93",X"00",X"00",X"00",X"00",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"ad",X"ad",X"ad",X"93",X"93",X"00",X"00",X"00",X"00",
    X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"ad",X"ad",X"ad",X"ad",X"00",X"00",X"00",X"00",X"00",
    X"16",X"5b",X"16",X"93",X"93",X"16",X"5b",X"ad",X"45",X"45",X"45",X"00",X"00",X"00",X"00",X"00",
    X"16",X"16",X"45",X"e5",X"93",X"16",X"5b",X"ad",X"93",X"16",X"16",X"5b",X"00",X"00",X"00",X"00",
    X"16",X"45",X"45",X"45",X"45",X"16",X"5b",X"ad",X"93",X"16",X"16",X"93",X"00",X"00",X"00",X"00",
    X"16",X"45",X"45",X"45",X"45",X"45",X"5b",X"ad",X"93",X"83",X"83",X"5b",X"00",X"00",X"00",X"00",
    X"16",X"45",X"45",X"45",X"45",X"45",X"5b",X"ad",X"93",X"e5",X"e5",X"00",X"00",X"00",X"00",X"00",
    X"16",X"45",X"45",X"45",X"16",X"45",X"5b",X"ad",X"93",X"16",X"16",X"00",X"00",X"00",X"00",X"00",
    X"16",X"45",X"16",X"45",X"45",X"45",X"5b",X"ad",X"93",X"93",X"93",X"00",X"00",X"00",X"00",X"00",
    X"16",X"93",X"93",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"93",X"93",X"16",X"16",
    X"93",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"93",X"93",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"45",X"ad",X"ad",X"ad",X"16",X"16",X"16",X"16",X"ad",X"5b",X"5b",X"45",X"45",X"45",X"16",X"16",
    X"ad",X"45",X"45",X"ad",X"93",X"93",X"93",X"93",X"ad",X"5b",X"5b",X"5b",X"45",X"45",X"16",X"16",
    X"45",X"93",X"16",X"45",X"ad",X"93",X"93",X"93",X"83",X"5b",X"5b",X"5b",X"45",X"45",X"16",X"16",
    X"00",X"93",X"16",X"16",X"45",X"ad",X"ad",X"ad",X"83",X"5b",X"5b",X"45",X"45",X"45",X"45",X"16",
    X"00",X"00",X"93",X"16",X"45",X"ad",X"ad",X"16",X"83",X"5b",X"5b",X"45",X"16",X"16",X"45",X"16",
    X"00",X"00",X"93",X"16",X"16",X"45",X"ad",X"93",X"83",X"5b",X"5b",X"16",X"45",X"45",X"45",X"16",
    X"00",X"00",X"00",X"93",X"16",X"45",X"ad",X"93",X"83",X"5b",X"5b",X"16",X"16",X"16",X"16",X"16",
    X"00",X"00",X"00",X"93",X"93",X"ad",X"ad",X"ad",X"ad",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"00",X"00",X"00",X"00",X"ad",X"ad",X"ad",X"ad",X"ad",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",
    X"00",X"00",X"00",X"00",X"45",X"45",X"45",X"ad",X"ad",X"5b",X"16",X"16",X"16",X"16",X"5b",X"16",
    X"00",X"00",X"00",X"5b",X"93",X"16",X"45",X"ad",X"ad",X"5b",X"16",X"16",X"16",X"45",X"16",X"16",
    X"00",X"00",X"00",X"93",X"93",X"16",X"45",X"ad",X"ad",X"5b",X"16",X"45",X"16",X"45",X"45",X"16",
    X"00",X"00",X"00",X"5b",X"93",X"16",X"45",X"ad",X"ad",X"5b",X"45",X"45",X"45",X"45",X"45",X"16",
    X"00",X"00",X"00",X"00",X"93",X"16",X"45",X"ad",X"ad",X"5b",X"45",X"45",X"45",X"45",X"45",X"16",
    X"00",X"00",X"00",X"00",X"93",X"16",X"45",X"ad",X"ad",X"5b",X"45",X"45",X"45",X"45",X"45",X"16",
    X"00",X"00",X"00",X"00",X"93",X"93",X"93",X"ad",X"ad",X"5b",X"45",X"45",X"45",X"45",X"45",X"16",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"2e",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"19",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"7b",X"2e",X"7b",X"19",X"19",X"19",X"19",X"19",X"4d",X"7b",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"7b",X"7b",X"2e",X"7b",X"19",X"19",X"19",X"19",X"19",X"7b",
    X"16",X"5b",X"5b",X"e5",X"e5",X"16",X"7b",X"2e",X"7b",X"19",X"7b",X"19",X"19",X"7b",X"19",X"19",
    X"16",X"e5",X"5b",X"e5",X"e5",X"16",X"2e",X"7b",X"7b",X"19",X"2e",X"19",X"2e",X"7b",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"2e",X"7b",X"2e",X"19",X"7b",X"19",X"2e",X"7b",X"19",X"19",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"19",X"19",X"7b",X"4d",X"4d",X"19",X"4d",X"7b",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"7b",X"4d",X"19",X"4d",X"19",X"19",X"4d",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"e5",X"e5",X"16",X"7b",X"19",X"19",X"7b",X"19",X"19",X"4d",X"19",X"19",X"19",
    X"16",X"e5",X"e5",X"5b",X"e5",X"16",X"7b",X"4d",X"19",X"19",X"19",X"7b",X"19",X"19",X"19",X"19",
    X"16",X"e5",X"5b",X"e5",X"5b",X"16",X"4d",X"2e",X"19",X"19",X"19",X"7b",X"4d",X"19",X"4d",X"19",
    X"16",X"e5",X"e5",X"5b",X"5b",X"16",X"7b",X"7b",X"19",X"4d",X"19",X"19",X"7b",X"19",X"19",X"4d",
    X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",X"4d",X"4d",X"4d",X"4d",X"19",X"4d",X"19",X"19",X"7b",
    X"16",X"45",X"16",X"83",X"83",X"16",X"45",X"16",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"19",
    X"19",X"4d",X"19",X"19",X"00",X"45",X"e5",X"5b",X"16",X"5b",X"e5",X"5b",X"00",X"19",X"19",X"19",
    X"19",X"4d",X"19",X"19",X"83",X"83",X"16",X"16",X"83",X"16",X"16",X"93",X"83",X"19",X"19",X"19",
    X"19",X"4d",X"4d",X"19",X"19",X"83",X"83",X"19",X"2e",X"19",X"83",X"83",X"19",X"19",X"7b",X"19",
    X"19",X"19",X"4d",X"19",X"19",X"00",X"00",X"2e",X"7b",X"4d",X"00",X"00",X"2e",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"7b",X"00",X"2e",X"7b",X"2e",X"00",X"19",X"4d",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"7b",X"19",X"7b",X"2e",X"2e",X"19",X"2e",X"2e",X"7b",X"7b",X"7b",
    X"2e",X"19",X"7b",X"19",X"19",X"2e",X"19",X"7b",X"2e",X"2e",X"2e",X"7b",X"2e",X"19",X"2e",X"2e",
    X"2e",X"19",X"7b",X"7b",X"19",X"2e",X"7b",X"2e",X"2e",X"2e",X"7b",X"7b",X"19",X"19",X"2e",X"19",
    X"2e",X"19",X"19",X"4d",X"2e",X"2e",X"2e",X"2e",X"4d",X"2e",X"2e",X"2e",X"19",X"2e",X"2e",X"19",
    X"4d",X"2e",X"19",X"7b",X"4d",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"7b",X"7b",X"19",X"19",X"19",
    X"4d",X"19",X"19",X"7b",X"7b",X"19",X"2e",X"19",X"2e",X"7b",X"2e",X"19",X"2e",X"19",X"19",X"4d",
    X"19",X"19",X"7b",X"19",X"4d",X"19",X"7b",X"4d",X"7b",X"19",X"19",X"2e",X"7b",X"19",X"4d",X"4d",
    X"19",X"19",X"2e",X"19",X"7b",X"19",X"7b",X"2e",X"19",X"19",X"2e",X"2e",X"4d",X"2e",X"4d",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"7b",X"19",X"19",X"19",X"2e",X"4d",X"19",X"2e",
    X"4d",X"19",X"19",X"19",X"4d",X"7b",X"7b",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"7b",X"7b",X"19",X"19",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"19",X"19",X"7b",
    X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"19",X"2e",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"4d",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"19",X"7b",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"19",X"19",X"19",X"4d",X"19",X"19",X"4d",X"19",X"19",X"4d",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"19",X"4d",X"4d",X"19",X"4d",X"19",X"4d",X"19",X"19",X"19",X"16",X"e5",X"e5",X"5b",X"5b",X"16",
    X"19",X"19",X"2e",X"19",X"4d",X"19",X"19",X"19",X"19",X"19",X"16",X"e5",X"e5",X"5b",X"e5",X"16",
    X"7b",X"19",X"2e",X"19",X"4d",X"19",X"19",X"19",X"19",X"4d",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"19",X"2e",X"4d",X"19",X"4d",X"19",X"19",X"19",X"7b",X"19",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"19",X"7b",X"4d",X"19",X"19",X"19",X"19",X"19",X"7b",X"7b",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"19",X"19",X"4d",X"19",X"19",X"4d",X"19",X"19",X"4d",X"2e",X"16",X"e5",X"e5",X"e5",X"e5",X"16",
    X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"7b",X"2e",X"16",X"e5",X"5b",X"e5",X"e5",X"16",
    X"19",X"19",X"19",X"19",X"19",X"4d",X"19",X"19",X"7b",X"2e",X"16",X"5b",X"e5",X"5b",X"e5",X"16",
    X"4d",X"19",X"19",X"19",X"4d",X"4d",X"19",X"19",X"4d",X"7b",X"16",X"5b",X"5b",X"e5",X"e5",X"16",
    X"4d",X"4d",X"19",X"2e",X"4d",X"19",X"4d",X"4d",X"4d",X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",
    X"7b",X"7b",X"19",X"19",X"19",X"19",X"19",X"2e",X"16",X"45",X"16",X"83",X"83",X"16",X"45",X"16",
    X"45",X"e5",X"5b",X"e5",X"e5",X"16",X"93",X"45",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"e5",X"16",
    X"45",X"e5",X"e5",X"e5",X"e5",X"16",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"45",X"e5",X"e5",X"e5",X"e5",X"16",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"45",X"e5",X"e5",X"5b",X"e5",X"16",X"93",X"45",X"16",X"00",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"45",X"e5",X"e5",X"5b",X"e5",X"16",X"93",X"16",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"45",X"5b",X"5b",X"e5",X"e5",X"16",X"93",X"5b",X"5b",X"83",X"45",X"5b",X"5b",X"e5",X"e5",X"16",
    X"45",X"e5",X"5b",X"e5",X"e5",X"16",X"93",X"45",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"e5",X"16",
    X"45",X"e5",X"e5",X"e5",X"e5",X"16",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"45",X"e5",X"e5",X"5b",X"e5",X"16",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"45",X"e5",X"e5",X"e5",X"e5",X"16",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"45",X"e5",X"e5",X"e5",X"e5",X"16",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"45",X"e5",X"e5",X"5b",X"e5",X"16",X"93",X"45",X"16",X"00",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"45",X"e5",X"5b",X"e5",X"5b",X"16",X"93",X"16",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"5b",X"16",
    X"45",X"e5",X"e5",X"5b",X"5b",X"16",X"93",X"5b",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"5b",X"16",
    X"45",X"e5",X"e5",X"e5",X"e5",X"16",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"45",X"e5",X"5b",X"e5",X"e5",X"16",X"93",X"45",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"e5",X"16",
    X"83",X"93",X"93",X"93",X"93",X"93",X"5b",X"5b",X"93",X"16",X"16",X"93",X"83",X"83",X"83",X"00",
    X"83",X"45",X"5b",X"93",X"e5",X"e5",X"45",X"45",X"93",X"16",X"16",X"83",X"16",X"83",X"00",X"83",
    X"83",X"16",X"45",X"93",X"5b",X"5b",X"45",X"45",X"93",X"93",X"93",X"83",X"93",X"83",X"00",X"83",
    X"83",X"16",X"45",X"93",X"5b",X"5b",X"93",X"93",X"93",X"45",X"45",X"83",X"93",X"00",X"83",X"83",
    X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"5b",X"5b",X"16",X"16",X"83",X"83",X"00",X"83",X"00",
    X"83",X"45",X"5b",X"e5",X"e5",X"e5",X"93",X"45",X"45",X"16",X"16",X"83",X"16",X"00",X"00",X"83",
    X"83",X"16",X"45",X"5b",X"5b",X"5b",X"93",X"45",X"45",X"93",X"93",X"16",X"93",X"00",X"00",X"83",
    X"83",X"16",X"45",X"5b",X"5b",X"5b",X"93",X"93",X"93",X"45",X"45",X"93",X"93",X"00",X"83",X"83",
    X"83",X"93",X"93",X"93",X"93",X"93",X"5b",X"5b",X"93",X"16",X"16",X"93",X"83",X"83",X"83",X"00",
    X"83",X"45",X"45",X"93",X"e5",X"e5",X"45",X"45",X"93",X"16",X"16",X"83",X"16",X"83",X"00",X"83",
    X"83",X"16",X"45",X"93",X"5b",X"5b",X"45",X"45",X"93",X"93",X"93",X"83",X"93",X"83",X"00",X"83",
    X"83",X"16",X"45",X"93",X"5b",X"5b",X"93",X"93",X"93",X"45",X"45",X"83",X"93",X"00",X"83",X"83",
    X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"5b",X"5b",X"16",X"16",X"83",X"83",X"00",X"83",X"00",
    X"83",X"45",X"5b",X"e5",X"e5",X"e5",X"93",X"45",X"45",X"16",X"16",X"83",X"16",X"00",X"00",X"83",
    X"83",X"16",X"45",X"5b",X"5b",X"5b",X"93",X"45",X"45",X"93",X"93",X"16",X"93",X"00",X"00",X"83",
    X"83",X"16",X"45",X"5b",X"5b",X"5b",X"93",X"93",X"93",X"45",X"45",X"93",X"93",X"00",X"83",X"83",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"4d",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"83",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"83",
    X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",
    X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",
    X"4d",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"16",X"16",X"16",X"83",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"83",X"16",X"16",X"16",X"16",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"4d",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",
    X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",
    X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",
    X"4d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"93",X"93",X"93",X"00",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"00",X"93",X"93",X"93",X"93",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"83",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"83",
    X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",
    X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"16",X"16",X"16",X"83",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"83",X"16",X"16",X"16",X"16",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",
    X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",
    X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"93",X"93",X"93",X"00",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"00",X"93",X"93",X"93",X"93",
    X"93",X"93",X"83",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5b",X"93",X"93",X"93",X"93",
    X"93",X"93",X"83",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5b",X"93",X"93",X"93",X"93",
    X"83",X"83",X"83",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5b",X"83",X"83",X"83",X"83",
    X"16",X"16",X"83",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5b",X"16",X"16",X"16",X"83",
    X"93",X"93",X"83",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5b",X"93",X"93",X"16",X"83",
    X"93",X"93",X"83",X"45",X"93",X"93",X"93",X"93",X"93",X"93",X"00",X"5b",X"93",X"93",X"16",X"83",
    X"83",X"83",X"83",X"45",X"93",X"16",X"16",X"16",X"16",X"16",X"83",X"5b",X"83",X"83",X"83",X"83",
    X"16",X"16",X"83",X"45",X"16",X"e5",X"e5",X"e5",X"e5",X"e5",X"83",X"5b",X"83",X"16",X"16",X"16",
    X"93",X"93",X"83",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"83",X"93",X"93",X"93",
    X"93",X"93",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",X"93",X"93",X"93",
    X"83",X"83",X"83",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"83",X"83",X"83",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",
    X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",
    X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"93",X"93",X"93",X"00",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"00",X"93",X"93",X"93",X"93",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"4d",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"83",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"4d",
    X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"4d",
    X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"4d",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"4d",
    X"16",X"16",X"16",X"83",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"83",X"16",X"16",X"16",X"16",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"93",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"4d",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"4d",
    X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"4d",
    X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"93",X"4d",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4d",
    X"93",X"93",X"93",X"00",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"00",X"93",X"93",X"93",X"93",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"93",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"45",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"16",X"45",X"93",X"45",X"16",X"83",X"83",X"93",X"83",
    X"16",X"5b",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"16",X"93",X"45",X"16",X"83",X"16",X"83",X"83",
    X"16",X"5b",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"5b",X"93",X"45",X"16",X"83",X"16",X"16",X"83",
    X"16",X"e5",X"e5",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"e5",X"5b",X"e5",X"45",X"83",X"5b",X"45",X"93",X"93",X"93",X"83",X"16",X"93",X"83",
    X"16",X"e5",X"5b",X"e5",X"e5",X"45",X"83",X"5b",X"45",X"93",X"45",X"93",X"83",X"16",X"93",X"83",
    X"16",X"16",X"16",X"16",X"16",X"45",X"83",X"5b",X"45",X"93",X"45",X"45",X"83",X"16",X"93",X"83",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"45",X"83",X"5b",X"45",X"93",X"45",X"16",X"83",X"16",X"93",X"83",
    X"5b",X"5b",X"e5",X"2e",X"2e",X"45",X"83",X"16",X"16",X"93",X"45",X"16",X"83",X"83",X"93",X"83",
    X"5b",X"5b",X"5b",X"5b",X"2e",X"45",X"83",X"5b",X"45",X"45",X"45",X"16",X"83",X"16",X"83",X"83",
    X"45",X"45",X"45",X"45",X"2e",X"45",X"83",X"45",X"e5",X"e5",X"2e",X"45",X"83",X"16",X"16",X"83",
    X"93",X"93",X"93",X"93",X"93",X"45",X"83",X"45",X"e5",X"e5",X"5b",X"2e",X"45",X"16",X"93",X"83",
    X"83",X"83",X"83",X"83",X"93",X"45",X"83",X"83",X"45",X"e5",X"e5",X"e5",X"2e",X"45",X"93",X"83",
    X"83",X"93",X"16",X"83",X"93",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"45",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"93",X"83",X"83",X"16",X"45",X"93",X"45",X"16",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"83",X"83",X"16",X"83",X"16",X"45",X"93",X"16",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"5b",X"16",
    X"83",X"16",X"16",X"83",X"16",X"45",X"93",X"5b",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"5b",X"16",
    X"83",X"93",X"16",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"93",X"93",X"93",X"45",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"93",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"45",X"45",X"93",X"45",X"5b",X"83",X"45",X"16",X"16",X"16",X"16",X"16",
    X"83",X"93",X"16",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"83",X"93",X"83",X"83",X"16",X"45",X"93",X"16",X"16",X"83",X"45",X"2e",X"2e",X"e5",X"5b",X"5b",
    X"83",X"83",X"16",X"83",X"16",X"45",X"45",X"45",X"5b",X"83",X"45",X"2e",X"5b",X"5b",X"5b",X"5b",
    X"83",X"16",X"16",X"83",X"45",X"2e",X"e5",X"e5",X"45",X"83",X"45",X"2e",X"45",X"45",X"45",X"45",
    X"83",X"93",X"16",X"45",X"2e",X"5b",X"e5",X"e5",X"45",X"83",X"45",X"93",X"93",X"93",X"93",X"93",
    X"83",X"93",X"45",X"2e",X"e5",X"e5",X"e5",X"45",X"83",X"83",X"45",X"93",X"83",X"83",X"83",X"83",
    X"16",X"45",X"45",X"45",X"45",X"45",X"5b",X"ad",X"ad",X"ad",X"ad",X"00",X"00",X"00",X"00",X"00",
    X"16",X"45",X"45",X"45",X"45",X"45",X"5b",X"ad",X"45",X"45",X"45",X"00",X"00",X"00",X"00",X"00",
    X"16",X"45",X"45",X"45",X"45",X"16",X"5b",X"ad",X"93",X"16",X"16",X"00",X"00",X"00",X"00",X"00",
    X"16",X"16",X"16",X"16",X"16",X"16",X"5b",X"ad",X"93",X"16",X"16",X"00",X"00",X"00",X"00",X"00",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"ad",X"93",X"16",X"16",X"00",X"00",X"00",X"00",X"00",
    X"16",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"ad",X"93",X"16",X"16",X"00",X"00",X"00",X"00",X"00",
    X"16",X"5b",X"16",X"16",X"16",X"16",X"5b",X"ad",X"93",X"16",X"16",X"00",X"00",X"00",X"00",X"00",
    X"16",X"16",X"16",X"45",X"45",X"16",X"5b",X"ad",X"93",X"93",X"93",X"00",X"00",X"00",X"00",X"00",
    X"16",X"45",X"45",X"45",X"45",X"45",X"5b",X"ad",X"ad",X"ad",X"ad",X"00",X"00",X"00",X"00",X"00",
    X"16",X"45",X"45",X"16",X"45",X"16",X"5b",X"ad",X"45",X"45",X"45",X"00",X"00",X"00",X"00",X"83",
    X"16",X"16",X"45",X"16",X"16",X"16",X"45",X"ad",X"93",X"16",X"16",X"00",X"00",X"00",X"00",X"83",
    X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"ad",X"93",X"16",X"16",X"5b",X"00",X"00",X"0a",X"0a",
    X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"ad",X"93",X"16",X"16",X"93",X"00",X"00",X"0a",X"0a",
    X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"ad",X"93",X"16",X"16",X"5b",X"00",X"0a",X"0a",X"0a",
    X"93",X"16",X"16",X"16",X"16",X"16",X"93",X"ad",X"93",X"16",X"16",X"00",X"0a",X"0a",X"0f",X"0f",
    X"93",X"93",X"93",X"93",X"93",X"93",X"ad",X"0a",X"ad",X"93",X"93",X"00",X"0a",X"0a",X"0f",X"0a",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"0a",X"83",X"0a",X"0a",X"0a",X"0a",X"0a",X"83",X"83",X"0a",X"0a",X"0a",X"0a",X"0a",X"83",X"0a",
    X"0a",X"83",X"83",X"0a",X"83",X"83",X"83",X"0a",X"0a",X"83",X"83",X"83",X"0a",X"83",X"83",X"0a",
    X"0a",X"0a",X"83",X"83",X"83",X"0a",X"83",X"0a",X"0a",X"83",X"0a",X"83",X"83",X"83",X"0a",X"0a",
    X"0a",X"0f",X"0f",X"0a",X"0a",X"0a",X"0a",X"0f",X"0f",X"0a",X"0a",X"0a",X"0a",X"0f",X"0f",X"0a",
    X"0a",X"0a",X"0f",X"0f",X"0a",X"0a",X"0f",X"0f",X"0f",X"0f",X"0a",X"0a",X"0f",X"0f",X"0a",X"0a",
    X"0a",X"0a",X"0a",X"0f",X"0f",X"0a",X"0a",X"0f",X"0f",X"0a",X"0a",X"0f",X"0f",X"0a",X"0a",X"0a",
    X"0f",X"0f",X"0a",X"0a",X"0f",X"0f",X"0a",X"0a",X"0a",X"0a",X"0f",X"0f",X"0a",X"0a",X"0f",X"0f",
    X"0a",X"0f",X"0a",X"0a",X"0a",X"0f",X"0f",X"0f",X"0f",X"0f",X"0f",X"0a",X"0a",X"0a",X"0f",X"0a",
    X"00",X"00",X"00",X"00",X"ad",X"ad",X"ad",X"ad",X"ad",X"5b",X"45",X"45",X"45",X"45",X"45",X"16",
    X"00",X"00",X"00",X"00",X"45",X"45",X"45",X"ad",X"ad",X"5b",X"16",X"45",X"45",X"45",X"45",X"16",
    X"00",X"00",X"00",X"00",X"93",X"16",X"45",X"ad",X"ad",X"5b",X"16",X"45",X"16",X"45",X"16",X"16",
    X"00",X"00",X"00",X"00",X"93",X"16",X"45",X"ad",X"ad",X"5b",X"16",X"16",X"16",X"16",X"16",X"16",
    X"00",X"00",X"00",X"00",X"93",X"16",X"45",X"ad",X"ad",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
    X"00",X"00",X"00",X"00",X"93",X"16",X"45",X"ad",X"ad",X"5b",X"5b",X"5b",X"5b",X"5b",X"5b",X"16",
    X"00",X"00",X"00",X"00",X"93",X"16",X"45",X"ad",X"ad",X"5b",X"16",X"16",X"16",X"16",X"16",X"16",
    X"00",X"00",X"00",X"00",X"93",X"93",X"93",X"ad",X"ad",X"5b",X"16",X"45",X"45",X"45",X"45",X"16",
    X"00",X"00",X"00",X"00",X"ad",X"ad",X"ad",X"ad",X"ad",X"5b",X"45",X"45",X"45",X"45",X"45",X"16",
    X"00",X"00",X"00",X"00",X"45",X"45",X"45",X"ad",X"ad",X"5b",X"16",X"45",X"16",X"45",X"45",X"16",
    X"00",X"00",X"00",X"00",X"93",X"16",X"45",X"ad",X"ad",X"45",X"16",X"16",X"16",X"45",X"16",X"16",
    X"0a",X"00",X"00",X"5b",X"93",X"16",X"45",X"ad",X"ad",X"45",X"16",X"16",X"16",X"16",X"16",X"16",
    X"0a",X"00",X"00",X"93",X"93",X"16",X"45",X"ad",X"83",X"45",X"16",X"16",X"16",X"16",X"16",X"16",
    X"0a",X"0a",X"00",X"5b",X"93",X"16",X"45",X"ad",X"83",X"45",X"16",X"16",X"16",X"16",X"16",X"16",
    X"0f",X"0f",X"0a",X"00",X"93",X"16",X"45",X"ad",X"83",X"93",X"16",X"16",X"16",X"16",X"16",X"93",
    X"0a",X"0f",X"0a",X"00",X"93",X"93",X"93",X"ad",X"0a",X"0a",X"93",X"93",X"93",X"93",X"93",X"93",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",
    X"45",X"5b",X"5b",X"e5",X"45",X"5b",X"e5",X"e5",X"45",X"2e",X"5b",X"e5",X"e5",X"e5",X"e5",X"16",
    X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",X"e5",X"5b",X"e5",X"45",X"2e",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"93",X"45",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"93",X"5b",X"83",X"45",X"e5",X"16",X"2e",X"e5",X"16",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"45",X"5b",X"83",X"45",X"e5",X"16",X"2e",X"e5",X"16",
    X"16",X"16",X"16",X"83",X"16",X"16",X"83",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"93",X"93",X"16",X"83",X"93",X"45",X"83",X"45",X"83",X"83",X"45",X"93",X"e5",X"5b",X"e5",X"16",
    X"83",X"83",X"83",X"83",X"16",X"45",X"83",X"83",X"5b",X"83",X"2e",X"2e",X"e5",X"5b",X"e5",X"16",
    X"93",X"93",X"83",X"83",X"16",X"45",X"83",X"5b",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"83",X"16",X"83",X"16",X"45",X"83",X"45",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"e5",X"16",
    X"83",X"93",X"16",X"83",X"16",X"83",X"83",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"93",X"93",X"16",X"83",X"93",X"93",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"83",X"83",X"83",X"83",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"16",X"16",X"16",X"16",X"16",X"45",X"93",X"45",X"16",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"93",X"93",X"93",X"93",X"16",X"45",X"93",X"16",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"5b",X"16",
    X"93",X"93",X"93",X"93",X"16",X"45",X"93",X"5b",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"5b",X"16",
    X"83",X"83",X"83",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"16",X"16",X"16",X"83",X"16",X"83",X"93",X"45",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"e5",X"16",
    X"93",X"93",X"16",X"83",X"83",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"93",X"93",X"83",X"83",X"45",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"83",X"83",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"93",X"83",X"16",X"83",X"16",X"45",X"93",X"45",X"16",X"83",X"45",X"e5",X"e5",X"5b",X"e5",X"16",
    X"83",X"83",X"16",X"83",X"16",X"45",X"93",X"16",X"5b",X"83",X"45",X"e5",X"5b",X"5b",X"e5",X"16",
    X"83",X"83",X"16",X"83",X"16",X"45",X"93",X"5b",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"e5",X"16",
    X"00",X"93",X"16",X"83",X"16",X"45",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"00",X"93",X"16",X"83",X"16",X"83",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",
    X"45",X"5b",X"5b",X"e5",X"45",X"5b",X"e5",X"e5",X"45",X"2e",X"5b",X"e5",X"e5",X"e5",X"e5",X"16",
    X"e5",X"e5",X"e5",X"5b",X"e5",X"e5",X"5b",X"e5",X"e5",X"e5",X"e5",X"5b",X"e5",X"45",X"2e",X"16",
    X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"e5",X"16",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"5b",X"5b",X"5b",X"5b",X"83",X"5b",X"5b",X"5b",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"45",X"45",X"45",X"45",X"16",X"5b",X"45",X"45",X"45",X"83",X"45",X"e5",X"16",X"2e",X"e5",X"16",
    X"16",X"16",X"16",X"16",X"93",X"5b",X"16",X"16",X"16",X"83",X"45",X"e5",X"16",X"2e",X"e5",X"16",
    X"93",X"93",X"93",X"93",X"83",X"93",X"93",X"93",X"93",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"5b",X"5b",X"83",X"93",X"93",X"e5",X"5b",X"e5",X"16",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"5b",X"83",X"2e",X"2e",X"e5",X"5b",X"e5",X"16",
    X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"45",X"5b",X"83",X"45",X"e5",X"5b",X"e5",X"e5",X"16",
    X"16",X"16",X"16",X"93",X"16",X"16",X"93",X"45",X"5b",X"83",X"45",X"e5",X"e5",X"e5",X"e5",X"16",
    X"83",X"93",X"93",X"93",X"93",X"93",X"5b",X"5b",X"93",X"16",X"16",X"93",X"83",X"83",X"83",X"19",
    X"83",X"45",X"45",X"93",X"e5",X"e5",X"45",X"45",X"93",X"16",X"16",X"83",X"16",X"83",X"83",X"7b",
    X"83",X"16",X"45",X"93",X"5b",X"5b",X"45",X"45",X"93",X"93",X"93",X"83",X"93",X"83",X"2e",X"7b",
    X"83",X"16",X"45",X"93",X"5b",X"5b",X"93",X"93",X"93",X"45",X"45",X"83",X"93",X"2e",X"7b",X"19",
    X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"5b",X"5b",X"16",X"16",X"83",X"2e",X"7b",X"19",X"19",
    X"83",X"45",X"45",X"e5",X"e5",X"e5",X"93",X"45",X"45",X"16",X"16",X"7b",X"19",X"19",X"19",X"19",
    X"83",X"16",X"45",X"5b",X"5b",X"5b",X"7b",X"45",X"45",X"2e",X"7b",X"4d",X"19",X"19",X"19",X"19",
    X"83",X"16",X"45",X"5b",X"5b",X"5b",X"7b",X"7b",X"2e",X"7b",X"19",X"4d",X"19",X"19",X"19",X"19",
    X"2e",X"2e",X"7b",X"7b",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"7b",X"19",X"19",
    X"7b",X"7b",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"4d",X"7b",X"19",X"19",X"19",X"19",
    X"19",X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"7b",X"7b",X"7b",X"7b",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"7b",X"7b",X"7b",X"7b",X"7b",X"19",X"19",X"19",X"4d",X"4d",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",
    X"4d",X"4d",X"19",X"4d",X"4d",X"7b",X"7b",X"19",X"7b",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",
    X"7b",X"7b",X"19",X"7b",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"83",X"93",X"93",X"93",X"93",X"93",X"5b",X"5b",X"93",X"16",X"16",X"93",X"83",X"83",X"83",X"19",
    X"83",X"45",X"45",X"93",X"e5",X"e5",X"45",X"45",X"93",X"16",X"16",X"83",X"16",X"83",X"83",X"4d",
    X"83",X"16",X"45",X"93",X"5b",X"5b",X"45",X"45",X"93",X"93",X"93",X"83",X"93",X"83",X"7b",X"19",
    X"83",X"16",X"45",X"93",X"5b",X"5b",X"93",X"93",X"93",X"45",X"45",X"83",X"93",X"2e",X"4d",X"19",
    X"83",X"93",X"93",X"93",X"93",X"93",X"93",X"5b",X"5b",X"16",X"16",X"83",X"2e",X"7b",X"19",X"19",
    X"83",X"45",X"45",X"e5",X"e5",X"e5",X"93",X"45",X"45",X"16",X"16",X"7b",X"4d",X"19",X"19",X"19",
    X"83",X"16",X"45",X"5b",X"5b",X"5b",X"7b",X"45",X"45",X"2e",X"2e",X"19",X"4d",X"19",X"19",X"19",
    X"83",X"16",X"45",X"5b",X"5b",X"5b",X"7b",X"4d",X"4d",X"19",X"19",X"19",X"4d",X"19",X"19",X"19",
    X"19",X"19",X"4d",X"7b",X"2e",X"2e",X"2e",X"4d",X"4d",X"4d",X"4d",X"19",X"7b",X"19",X"19",X"19",
    X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"4d",X"7b",X"19",X"19",X"19",X"19",X"19",
    X"19",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"7b",X"7b",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",
    X"19",X"7b",X"7b",X"7b",X"7b",X"7b",X"19",X"19",X"19",X"19",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"19",X"19",X"19",X"19",X"19",X"19",X"4d",X"4d",X"19",X"4d",X"4d",X"4d",X"19",X"19",X"19",X"19",
    X"19",X"4d",X"4d",X"19",X"4d",X"4d",X"4d",X"4d",X"19",X"4d",X"4d",X"7b",X"19",X"19",X"19",X"19",
    X"19",X"4d",X"4d",X"19",X"4d",X"4d",X"7b",X"7b",X"19",X"7b",X"7b",X"19",X"19",X"19",X"19",X"19",
    X"19",X"7b",X"7b",X"19",X"7b",X"7b",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",    others=>X"01"
    );
end package;