use work.graphics_pkg.all;

package bomberman_pkg is
    constant BOMBERMAN_WIDTH : integer := 16;
    constant BOMBERMAN_HEIGHT : integer := 32;
    type bomberman_bitmap_type is array (0 to BOMBERMAN_HEIGHT-1, 0 to BOMBERMAN_WIDTH-1) of pixel_type;
    type bomberman_rom_type is array(0 to 2**14 -1) of pixel_type;
    
    constant BOMBERMAN_FRAMES : bomberman_rom_type :=
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"6a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"5a",X"5a",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"5a",X"5a",X"2e",X"5a",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"a5",X"21",X"21",X"a5",X"5a",X"5a",X"5a",X"5a",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"6a",X"a5",X"21",X"21",X"a5",X"a5",X"5a",X"5a",X"a5",X"21",X"21",X"21",X"a5",X"6a",X"01",
        X"01",X"6a",X"a5",X"a5",X"21",X"21",X"a5",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",
        X"01",X"6a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01",X"01",
        X"01",X"01",X"6a",X"6a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"a5",X"6a",X"6a",X"01",X"01",X"01",
        X"01",X"6a",X"9a",X"00",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"b2",X"c7",X"6a",X"01",X"01",
        X"01",X"c7",X"9a",X"00",X"b2",X"b2",X"b2",X"d8",X"d8",X"2e",X"d8",X"b2",X"9a",X"9a",X"01",X"01",
        X"01",X"5a",X"5a",X"00",X"b2",X"b2",X"d8",X"d8",X"d8",X"d8",X"d8",X"00",X"5a",X"5a",X"01",X"01",
        X"01",X"5a",X"5a",X"b2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"b2",X"5a",X"5a",X"01",X"01",
        X"01",X"01",X"01",X"c7",X"b2",X"b2",X"b2",X"d8",X"d8",X"d8",X"b2",X"c7",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"9a",X"9a",X"b2",X"b2",X"b2",X"b2",X"b2",X"9a",X"9a",X"01",X"01",X"01",X"01",
        X"01",X"01",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"c7",X"9a",X"9a",X"00",X"01",X"01",X"01",
        X"01",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"5a",X"5a",X"a5",X"01",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"5a",X"5a",X"2e",X"5a",X"a5",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"5a",X"5a",X"5a",X"5a",X"a5",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"a5",X"5a",X"5a",X"a5",X"a5",X"01",
        X"6a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"a5",X"a5",X"a5",X"6a",X"01",
        X"6a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",
        X"01",X"6a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01",X"01",
        X"01",X"c7",X"6a",X"6a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"a5",X"a5",X"6a",X"01",X"01",X"01",
        X"01",X"9a",X"9a",X"00",X"00",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"c7",X"9a",X"6a",X"01",X"01",
        X"01",X"6a",X"9a",X"00",X"b2",X"b2",X"b2",X"d8",X"d8",X"2e",X"d8",X"9a",X"9a",X"9a",X"01",X"01",
        X"01",X"01",X"6a",X"00",X"b2",X"b2",X"d8",X"d8",X"d8",X"d8",X"d8",X"5a",X"2e",X"5a",X"01",X"01",
        X"01",X"01",X"01",X"b2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"01",X"01",
        X"01",X"01",X"01",X"c7",X"b2",X"b2",X"b2",X"d8",X"d8",X"d8",X"b2",X"5a",X"5a",X"5a",X"01",X"01",
        X"01",X"01",X"00",X"9a",X"9a",X"b2",X"b2",X"b2",X"d8",X"b2",X"c7",X"6a",X"01",X"01",X"01",X"01",
        X"01",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"01",X"01",X"01",
        X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"00",X"00",X"00",X"c7",X"9a",X"9a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"01",X"6a",X"5a",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",
        X"6a",X"5a",X"5a",X"2e",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"5a",X"5a",X"5a",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"5a",X"5a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"6a",X"a5",X"a5",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01",
        X"6a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",
        X"01",X"6a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01",X"01",
        X"01",X"01",X"6a",X"6a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"a5",X"a5",X"6a",X"9a",X"01",X"01",
        X"01",X"6a",X"9a",X"9a",X"00",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"b2",X"c7",X"9a",X"01",X"01",
        X"01",X"c7",X"9a",X"9a",X"b2",X"b2",X"b2",X"d8",X"d8",X"2e",X"d8",X"b2",X"9a",X"6a",X"01",X"01",
        X"01",X"5a",X"2e",X"5a",X"b2",X"b2",X"d8",X"d8",X"d8",X"d8",X"d8",X"00",X"6a",X"01",X"01",X"01",
        X"01",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"b2",X"01",X"01",X"01",X"01",
        X"01",X"5a",X"5a",X"5a",X"b2",X"b2",X"b2",X"d8",X"d8",X"d8",X"b2",X"c7",X"01",X"01",X"01",X"01",
        X"01",X"01",X"00",X"6a",X"c7",X"b2",X"b2",X"b2",X"d8",X"b2",X"9a",X"9a",X"01",X"01",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"c7",X"9a",X"9a",X"00",X"01",X"01",X"01",
        X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"5a",X"5a",X"2e",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"5a",X"5a",X"5a",X"5a",X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"5a",X"5a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"21",X"a5",
        X"01",X"01",X"6a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"4e",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"4e",X"31",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"31",X"00",X"31",X"01",
        X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"31",X"00",X"31",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"31",X"00",X"31",X"4e",
        X"01",X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"31",X"00",X"4e",X"01",
        X"01",X"01",X"01",X"6a",X"a5",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"4e",X"4e",X"6a",X"01",
        X"01",X"01",X"01",X"01",X"b2",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"01",X"01",
        X"01",X"01",X"01",X"01",X"b2",X"d8",X"b2",X"c7",X"9a",X"9a",X"b2",X"2e",X"b2",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"d8",X"b2",X"9a",X"9a",X"9a",X"d8",X"d8",X"31",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"b2",X"00",X"00",X"5a",X"2e",X"5a",X"00",X"00",X"b2",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"b2",X"b2",X"5a",X"5a",X"5a",X"d8",X"b2",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"00",X"00",X"00",X"b2",X"5a",X"5a",X"5a",X"b2",X"5a",X"00",X"01",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"5a",X"c7",X"9a",X"9a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"2e",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"5a",X"5a",X"2e",X"5a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01",
        X"5a",X"5a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"4e",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"4e",X"4e",X"01",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"4e",X"4e",X"4e",X"31",X"00",X"01",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"4e",X"31",X"31",X"00",X"31",X"31",X"00",X"01",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"4e",X"31",X"31",X"00",X"31",X"31",X"00",X"01",X"01",
        X"01",X"a5",X"a5",X"21",X"21",X"21",X"21",X"4e",X"31",X"31",X"00",X"31",X"31",X"00",X"4e",X"01",
        X"01",X"6a",X"a5",X"a5",X"a5",X"21",X"21",X"4e",X"31",X"31",X"00",X"31",X"4e",X"4e",X"01",X"01",
        X"01",X"01",X"6a",X"6a",X"a5",X"a5",X"a5",X"6a",X"4e",X"4e",X"4e",X"4e",X"6a",X"6a",X"01",X"01",
        X"01",X"01",X"5a",X"00",X"00",X"6a",X"6a",X"6a",X"6a",X"6a",X"5a",X"2e",X"5a",X"01",X"01",X"01",
        X"01",X"01",X"5a",X"b2",X"b2",X"d8",X"b2",X"c7",X"9a",X"9a",X"5a",X"5a",X"5a",X"01",X"01",X"01",
        X"01",X"01",X"01",X"00",X"b2",X"d8",X"b2",X"b2",X"9a",X"9a",X"5a",X"5a",X"5a",X"01",X"01",X"01",
        X"01",X"01",X"01",X"b2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"b2",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"00",X"b2",X"b2",X"9a",X"9a",X"d8",X"b2",X"b2",X"c7",X"00",X"01",X"01",X"01",
        X"01",X"01",X"00",X"00",X"5a",X"c7",X"9a",X"9a",X"6a",X"b2",X"6a",X"9a",X"9a",X"5a",X"5a",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"9a",X"9a",X"6a",X"00",X"00",X"6a",X"6a",X"5a",X"5a",X"5a",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"5a",X"6a",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"2e",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"00",X"00",X"00",
        X"01",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
        X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",
        X"01",X"5a",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"4e",
        X"5a",X"5a",X"2e",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",
        X"5a",X"5a",X"5a",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",
        X"01",X"5a",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"4e",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"4e",X"01",
        X"01",X"01",X"01",X"6a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"a5",X"6a",X"5a",X"5a",
        X"01",X"01",X"01",X"01",X"00",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"b2",X"6a",X"5a",X"5a",
        X"01",X"01",X"01",X"01",X"b2",X"00",X"b2",X"9a",X"9a",X"b2",X"2e",X"d8",X"b2",X"6a",X"5a",X"5a",
        X"01",X"01",X"01",X"01",X"b2",X"b2",X"c7",X"9a",X"b2",X"d8",X"d8",X"b2",X"31",X"01",X"01",X"01",
        X"01",X"01",X"00",X"6a",X"5a",X"2e",X"5a",X"9a",X"00",X"00",X"00",X"00",X"b2",X"00",X"01",X"01",
        X"01",X"00",X"6a",X"c7",X"5a",X"5a",X"5a",X"6a",X"b2",X"9a",X"c7",X"b2",X"00",X"00",X"00",X"01",
        X"00",X"00",X"5a",X"9a",X"5a",X"5a",X"5a",X"b2",X"6a",X"9a",X"9a",X"9a",X"6a",X"5a",X"5a",X"00",
        X"00",X"00",X"5a",X"5a",X"9a",X"00",X"00",X"00",X"00",X"6a",X"9a",X"9a",X"5a",X"2e",X"5a",X"00",
        X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"9a",X"5a",X"5a",X"5a",X"00",X"00",
        X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",
        X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"00",X"00",X"00",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"2e",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"6a",X"6a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"a5",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"21",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"6a",X"01",
        X"01",X"6a",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"a5",X"01",X"01",
        X"01",X"6a",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"6a",X"01",X"01",
        X"01",X"01",X"6a",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"6a",X"01",X"01",X"01",
        X"01",X"6a",X"9a",X"00",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"00",X"c7",X"6a",X"01",X"01",
        X"01",X"c7",X"9a",X"00",X"b2",X"b2",X"d8",X"d8",X"d8",X"2e",X"d8",X"b2",X"9a",X"9a",X"01",X"01",
        X"01",X"5a",X"5a",X"00",X"b2",X"d8",X"d8",X"d8",X"d8",X"d8",X"d8",X"00",X"5a",X"5a",X"01",X"01",
        X"01",X"5a",X"5a",X"b2",X"00",X"00",X"31",X"31",X"31",X"00",X"00",X"b2",X"5a",X"5a",X"01",X"01",
        X"01",X"01",X"01",X"c7",X"b2",X"b2",X"d8",X"d8",X"d8",X"d8",X"b2",X"c7",X"01",X"01",X"01",X"01",
        X"01",X"01",X"00",X"9a",X"9a",X"b2",X"b2",X"d8",X"d8",X"b2",X"9a",X"9a",X"00",X"01",X"01",X"01",
        X"01",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"c7",X"9a",X"9a",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"2e",X"00",X"00",X"00",X"5a",X"5a",X"2e",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"5a",X"5a",X"2e",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"5a",X"5a",X"5a",X"5a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01",
        X"01",X"5a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"a5",X"21",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"4e",X"a5",X"01",
        X"6a",X"a5",X"a5",X"21",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"4e",X"a5",X"01",
        X"6a",X"6a",X"a5",X"a5",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"4e",X"6a",X"01",
        X"01",X"6a",X"6a",X"a5",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"4e",X"6a",X"01",
        X"01",X"01",X"6a",X"6a",X"6a",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"6a",X"01",X"01",
        X"01",X"6a",X"9a",X"00",X"00",X"6a",X"6a",X"6a",X"6a",X"5a",X"2e",X"5a",X"c7",X"9a",X"01",X"01",
        X"01",X"c7",X"9a",X"00",X"b2",X"b2",X"d8",X"d8",X"b2",X"5a",X"5a",X"5a",X"9a",X"6a",X"01",X"01",
        X"01",X"5a",X"5a",X"00",X"b2",X"d8",X"d8",X"d8",X"b2",X"5a",X"5a",X"5a",X"6a",X"01",X"01",X"01",
        X"01",X"01",X"01",X"9a",X"00",X"00",X"31",X"31",X"31",X"00",X"00",X"6a",X"01",X"01",X"01",X"01",
        X"01",X"01",X"00",X"c7",X"9a",X"b2",X"d8",X"d8",X"d8",X"b2",X"9a",X"6a",X"00",X"01",X"01",X"01",
        X"01",X"00",X"00",X"9a",X"9a",X"9a",X"b2",X"d8",X"b2",X"c7",X"9a",X"5a",X"00",X"00",X"01",X"01",
        X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"5a",X"00",X"00",X"01",X"01",X"01",
        X"00",X"00",X"5a",X"5a",X"2e",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
        X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
        X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"2e",X"5a",X"01",
        X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"5a",X"5a",X"5a",X"5a",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"5a",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"01",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"01",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"4e",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"4e",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"4e",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"21",X"a5",X"6a",X"01",
        X"6a",X"4e",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"a5",X"6a",X"01",X"01",
        X"01",X"6a",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"6a",X"6a",X"6a",X"01",X"01",X"01",
        X"01",X"c7",X"9a",X"5a",X"2e",X"5a",X"6a",X"6a",X"6a",X"6a",X"b2",X"b2",X"c7",X"6a",X"01",X"01",
        X"01",X"6a",X"9a",X"5a",X"5a",X"5a",X"b2",X"b2",X"d8",X"2e",X"d8",X"b2",X"9a",X"9a",X"01",X"01",
        X"01",X"01",X"6a",X"5a",X"5a",X"5a",X"b2",X"b2",X"d8",X"d8",X"d8",X"00",X"5a",X"5a",X"01",X"01",
        X"01",X"01",X"01",X"6a",X"00",X"00",X"31",X"31",X"31",X"00",X"00",X"c7",X"01",X"01",X"01",X"01",
        X"01",X"01",X"00",X"6a",X"c7",X"b2",X"b2",X"d8",X"d8",X"b2",X"9a",X"9a",X"01",X"01",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"9a",X"9a",X"b2",X"b2",X"b2",X"c7",X"9a",X"9a",X"00",X"01",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"00",X"5a",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"2e",X"5a",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"2e",X"5a",
        X"01",X"01",X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"5a",X"5a",X"5a",X"5a",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"5a",X"5a",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",
        X"4e",X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"01",X"31",X"4e",X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"01",X"31",X"00",X"31",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"01",X"31",X"00",X"31",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01",
        X"4e",X"31",X"00",X"31",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",
        X"01",X"4e",X"00",X"31",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01",X"01",
        X"01",X"6a",X"4e",X"4e",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"6a",X"6a",X"01",X"01",X"01",
        X"01",X"01",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"b2",X"b2",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"b2",X"d8",X"b2",X"c7",X"9a",X"9a",X"b2",X"2e",X"d8",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"31",X"d8",X"b2",X"9a",X"9a",X"9a",X"d8",X"d8",X"00",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"b2",X"00",X"00",X"5a",X"2e",X"5a",X"00",X"00",X"b2",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"00",X"b2",X"b2",X"5a",X"5a",X"5a",X"d8",X"b2",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"00",X"00",X"5a",X"b2",X"5a",X"5a",X"5a",X"b2",X"00",X"00",X"01",X"01",X"01",X"01",
        X"01",X"00",X"00",X"00",X"5a",X"5a",X"c7",X"9a",X"9a",X"5a",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"00",X"00",X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"2e",X"5a",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"4e",X"a5",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"5a",X"5a",X"01",
        X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"5a",X"5a",X"2e",X"5a",
        X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"5a",X"5a",X"5a",X"5a",
        X"4e",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"5a",X"5a",X"01",
        X"01",X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01",
        X"01",X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",
        X"01",X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01",X"01",
        X"5a",X"5a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"a5",X"6a",X"01",X"01",X"01",
        X"5a",X"5a",X"6a",X"b2",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"b2",X"01",X"01",X"01",X"01",
        X"5a",X"5a",X"6a",X"b2",X"d8",X"b2",X"6a",X"c7",X"9a",X"b2",X"b2",X"d8",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"31",X"d8",X"b2",X"b2",X"6a",X"9a",X"9a",X"d8",X"d8",X"01",X"01",X"01",X"01",
        X"01",X"01",X"00",X"b2",X"00",X"00",X"00",X"00",X"9a",X"5a",X"2e",X"5a",X"6a",X"01",X"01",X"01",
        X"01",X"00",X"00",X"00",X"b2",X"9a",X"9a",X"b2",X"6a",X"5a",X"5a",X"5a",X"9a",X"6a",X"01",X"01",
        X"00",X"5a",X"5a",X"6a",X"c7",X"9a",X"9a",X"b2",X"b2",X"5a",X"5a",X"5a",X"9a",X"5a",X"00",X"01",
        X"00",X"5a",X"2e",X"5a",X"9a",X"9a",X"6a",X"00",X"00",X"00",X"00",X"9a",X"5a",X"5a",X"00",X"01",
        X"00",X"00",X"5a",X"5a",X"5a",X"9a",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",
        X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"00",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",
        X"01",X"01",X"01",X"01",X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"a5",X"5a",X"5a",X"2e",X"5a",
        X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"5a",X"5a",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",
        X"01",X"4e",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"01",X"01",X"4e",X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",
        X"01",X"01",X"00",X"31",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",
        X"01",X"01",X"00",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",
        X"01",X"01",X"00",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",
        X"01",X"4e",X"00",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"01",X"6a",X"4e",X"4e",X"31",X"00",X"31",X"31",X"4e",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01",
        X"01",X"01",X"6a",X"6a",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"21",X"a5",X"6a",X"6a",X"01",X"01",
        X"01",X"01",X"01",X"5a",X"2e",X"5a",X"6a",X"6a",X"6a",X"6a",X"6a",X"b2",X"b2",X"5a",X"01",X"01",
        X"01",X"01",X"01",X"5a",X"5a",X"5a",X"c7",X"9a",X"9a",X"b2",X"d8",X"2e",X"d8",X"5a",X"01",X"01",
        X"01",X"01",X"01",X"5a",X"5a",X"5a",X"9a",X"9a",X"b2",X"b2",X"d8",X"d8",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"b2",X"31",X"00",X"00",X"00",X"00",X"00",X"00",X"b2",X"01",X"01",X"01",
        X"01",X"01",X"00",X"00",X"9a",X"b2",X"b2",X"b2",X"d8",X"c7",X"9a",X"b2",X"00",X"01",X"01",X"01",
        X"01",X"5a",X"5a",X"c7",X"9a",X"6a",X"b2",X"b2",X"6a",X"9a",X"9a",X"9a",X"5a",X"00",X"01",X"01",
        X"01",X"5a",X"5a",X"5a",X"6a",X"6a",X"00",X"00",X"00",X"6a",X"9a",X"9a",X"5a",X"5a",X"00",X"01",
        X"01",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"6a",X"5a",X"5a",X"2e",X"00",X"01",
        X"00",X"00",X"00",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"01",
        X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"00",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"2e",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"6a",X"6a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"a5",X"01",
        X"6a",X"a5",X"21",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"2e",X"2e",X"2e",X"31",X"2e",X"2e",X"2e",X"31",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"2e",X"00",X"2e",X"31",X"2e",X"00",X"2e",X"31",X"4e",X"21",X"6a",X"01",
        X"5a",X"5a",X"4e",X"31",X"2e",X"2e",X"2e",X"31",X"2e",X"2e",X"2e",X"31",X"4e",X"5a",X"5a",X"01",
        X"5a",X"5a",X"4e",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"4e",X"5a",X"5a",X"01",
        X"5a",X"5a",X"6a",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"c7",X"5a",X"5a",X"01",
        X"6a",X"c7",X"9a",X"00",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"00",X"9a",X"9a",X"6a",X"01",
        X"01",X"6a",X"9a",X"00",X"b2",X"b2",X"d8",X"d8",X"d8",X"2e",X"d8",X"b2",X"9a",X"6a",X"01",X"01",
        X"01",X"01",X"6a",X"00",X"b2",X"d8",X"d8",X"d8",X"d8",X"d8",X"d8",X"00",X"6a",X"01",X"01",X"01",
        X"01",X"01",X"01",X"b2",X"00",X"00",X"31",X"31",X"31",X"00",X"00",X"b2",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"c7",X"b2",X"b2",X"d8",X"d8",X"d8",X"d8",X"b2",X"c7",X"01",X"01",X"01",X"01",
        X"01",X"01",X"00",X"9a",X"9a",X"b2",X"b2",X"d8",X"d8",X"b2",X"9a",X"9a",X"00",X"01",X"01",X"01",
        X"01",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"c7",X"9a",X"9a",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"2e",X"00",X"00",X"00",X"5a",X"5a",X"2e",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"5a",X"5a",X"2e",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"5a",X"5a",X"5a",X"5a",X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"5a",X"5a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"21",X"4e",
        X"01",X"01",X"6a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"4e",X"31",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"31",X"2e",X"2e",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"5a",X"5a",X"5a",X"31",X"2e",X"00",X"01",
        X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"6a",X"5a",X"5a",X"5a",X"31",X"2e",X"2e",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"6a",X"5a",X"5a",X"5a",X"31",X"31",X"31",X"4e",
        X"01",X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"6a",X"c7",X"9a",X"6a",X"31",X"31",X"4e",X"01",
        X"01",X"01",X"01",X"6a",X"a5",X"a5",X"a5",X"21",X"6a",X"9a",X"9a",X"6a",X"4e",X"4e",X"6a",X"01",
        X"01",X"01",X"01",X"01",X"b2",X"6a",X"6a",X"6a",X"c7",X"9a",X"9a",X"6a",X"6a",X"6a",X"01",X"01",
        X"01",X"01",X"01",X"01",X"b2",X"d8",X"b2",X"b2",X"9a",X"9a",X"6a",X"2e",X"b2",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"d8",X"b2",X"b2",X"b2",X"b2",X"d8",X"d8",X"31",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"b2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"b2",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"b2",X"b2",X"b2",X"b2",X"b2",X"d8",X"b2",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"00",X"00",X"00",X"b2",X"b2",X"9a",X"b2",X"b2",X"5a",X"00",X"01",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"5a",X"c7",X"9a",X"9a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"2e",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"2e",X"5a",
        X"01",X"01",X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"5a",X"5a",X"5a",X"5a",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"5a",X"5a",X"01",
        X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"01",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",
        X"01",X"31",X"4e",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"01",X"2e",X"2e",X"31",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"01",X"00",X"2e",X"31",X"5a",X"5a",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"01",X"2e",X"2e",X"31",X"5a",X"5a",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01",
        X"4e",X"31",X"31",X"31",X"5a",X"5a",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",
        X"01",X"4e",X"31",X"31",X"6a",X"c7",X"9a",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01",X"01",
        X"01",X"6a",X"4e",X"4e",X"6a",X"9a",X"9a",X"6a",X"21",X"21",X"a5",X"6a",X"6a",X"01",X"01",X"01",
        X"01",X"01",X"6a",X"6a",X"6a",X"9a",X"9a",X"9a",X"6a",X"6a",X"b2",X"b2",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"b2",X"b2",X"6a",X"9a",X"9a",X"b2",X"b2",X"2e",X"d8",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"31",X"b2",X"b2",X"b2",X"b2",X"d8",X"d8",X"d8",X"00",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"b2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"b2",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"00",X"b2",X"b2",X"b2",X"b2",X"b2",X"d8",X"b2",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"00",X"00",X"5a",X"b2",X"b2",X"9a",X"b2",X"b2",X"00",X"00",X"01",X"01",X"01",X"01",
        X"01",X"00",X"00",X"00",X"5a",X"5a",X"c7",X"9a",X"9a",X"5a",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"00",X"00",X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"2e",X"5a",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"2e",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"01",X"6a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"21",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"2e",X"2e",X"2e",X"31",X"2e",X"2e",X"2e",X"31",X"4e",X"a5",X"6a",X"01",
        X"6a",X"6a",X"4e",X"31",X"2e",X"00",X"2e",X"31",X"2e",X"00",X"2e",X"31",X"4e",X"a5",X"6a",X"01",
        X"5a",X"5a",X"5a",X"31",X"2e",X"2e",X"2e",X"31",X"2e",X"2e",X"2e",X"31",X"5a",X"5a",X"5a",X"01",
        X"5a",X"5a",X"5a",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"5a",X"5a",X"5a",X"01",
        X"5a",X"5a",X"c7",X"00",X"b2",X"b2",X"b2",X"b2",X"d8",X"d8",X"d8",X"00",X"c7",X"5a",X"5a",X"01",
        X"01",X"6a",X"6a",X"b2",X"00",X"b2",X"b2",X"d8",X"d8",X"d8",X"00",X"b2",X"6a",X"6a",X"01",X"01",
        X"01",X"01",X"01",X"6a",X"b2",X"00",X"31",X"31",X"31",X"00",X"b2",X"6a",X"01",X"01",X"01",X"01",
        X"01",X"00",X"00",X"9a",X"6a",X"b2",X"b2",X"b2",X"d8",X"b2",X"6a",X"9a",X"00",X"01",X"01",X"01",
        X"00",X"00",X"00",X"c7",X"9a",X"6a",X"00",X"00",X"00",X"6a",X"c7",X"9a",X"00",X"00",X"01",X"01",
        X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"00",X"00",X"5a",X"5a",X"2e",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"2e",X"5a",X"00",X"01",X"01",
        X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"01",X"01",
        X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"2e",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"6a",X"6a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"a5",X"01",
        X"6a",X"a5",X"21",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"2e",X"2e",X"2e",X"31",X"2e",X"2e",X"2e",X"31",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"2e",X"00",X"2e",X"31",X"2e",X"00",X"2e",X"31",X"4e",X"21",X"6a",X"01",
        X"01",X"6a",X"4e",X"31",X"2e",X"2e",X"2e",X"31",X"2e",X"2e",X"2e",X"31",X"4e",X"a5",X"01",X"01",
        X"5a",X"5a",X"5a",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"5a",X"5a",X"5a",X"01",
        X"5a",X"5a",X"5a",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"5a",X"5a",X"5a",X"01",
        X"5a",X"5a",X"5a",X"00",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"00",X"5a",X"5a",X"5a",X"01",
        X"01",X"c7",X"9a",X"00",X"b2",X"b2",X"d8",X"d8",X"d8",X"2e",X"d8",X"b2",X"c7",X"9a",X"01",X"01",
        X"01",X"01",X"6a",X"00",X"b2",X"d8",X"d8",X"d8",X"d8",X"d8",X"d8",X"00",X"6a",X"01",X"01",X"01",
        X"01",X"00",X"00",X"b2",X"00",X"00",X"31",X"31",X"31",X"00",X"00",X"b2",X"00",X"00",X"01",X"01",
        X"00",X"00",X"5a",X"5a",X"c7",X"b2",X"d8",X"d8",X"d8",X"b2",X"9a",X"5a",X"5a",X"00",X"00",X"01",
        X"00",X"5a",X"5a",X"5a",X"5a",X"9a",X"b2",X"b2",X"b2",X"c7",X"5a",X"5a",X"5a",X"5a",X"00",X"01",
        X"00",X"5a",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"5a",X"00",X"01",
        X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"2e",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"6a",X"6a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"a5",X"01",
        X"6a",X"a5",X"21",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"2e",X"2e",X"2e",X"31",X"2e",X"2e",X"2e",X"31",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"2e",X"00",X"2e",X"31",X"2e",X"00",X"2e",X"31",X"4e",X"21",X"6a",X"01",
        X"01",X"6a",X"4e",X"31",X"2e",X"2e",X"2e",X"31",X"2e",X"2e",X"2e",X"31",X"4e",X"a5",X"01",X"01",
        X"5a",X"5a",X"5a",X"31",X"31",X"2e",X"31",X"31",X"31",X"31",X"31",X"31",X"5a",X"5a",X"5a",X"01",
        X"5a",X"5a",X"5a",X"4e",X"2e",X"2e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"5a",X"5a",X"5a",X"01",
        X"5a",X"5a",X"5a",X"00",X"2e",X"2e",X"6a",X"6a",X"6a",X"6a",X"6a",X"00",X"5a",X"5a",X"5a",X"01",
        X"01",X"c7",X"9a",X"00",X"b2",X"b2",X"d8",X"d8",X"d8",X"2e",X"d8",X"b2",X"c7",X"9a",X"01",X"01",
        X"01",X"01",X"6a",X"00",X"b2",X"d8",X"d8",X"d8",X"d8",X"d8",X"d8",X"00",X"6a",X"01",X"01",X"01",
        X"01",X"00",X"00",X"b2",X"00",X"00",X"31",X"31",X"31",X"00",X"00",X"b2",X"00",X"00",X"01",X"01",
        X"00",X"00",X"5a",X"5a",X"c7",X"b2",X"d8",X"d8",X"d8",X"b2",X"9a",X"5a",X"5a",X"00",X"00",X"01",
        X"00",X"5a",X"5a",X"5a",X"5a",X"9a",X"b2",X"b2",X"b2",X"c7",X"5a",X"5a",X"5a",X"5a",X"00",X"01",
        X"00",X"5a",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"5a",X"00",X"01",
        X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"2e",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"6a",X"6a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"a5",X"01",
        X"6a",X"a5",X"21",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"2e",X"2e",X"2e",X"31",X"2e",X"2e",X"2e",X"31",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"2e",X"00",X"2e",X"31",X"2e",X"00",X"2e",X"31",X"4e",X"21",X"6a",X"01",
        X"01",X"6a",X"4e",X"31",X"2e",X"2e",X"2e",X"31",X"2e",X"2e",X"2e",X"31",X"4e",X"a5",X"01",X"01",
        X"5a",X"5a",X"5a",X"31",X"31",X"2e",X"31",X"31",X"31",X"31",X"31",X"31",X"5a",X"5a",X"5a",X"01",
        X"5a",X"5a",X"5a",X"4e",X"4e",X"2e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"5a",X"5a",X"5a",X"01",
        X"5a",X"5a",X"5a",X"00",X"6a",X"2e",X"6a",X"6a",X"6a",X"6a",X"6a",X"00",X"5a",X"5a",X"5a",X"01",
        X"01",X"c7",X"9a",X"00",X"2e",X"2e",X"d8",X"d8",X"d8",X"2e",X"d8",X"b2",X"c7",X"9a",X"01",X"01",
        X"01",X"01",X"6a",X"00",X"2e",X"2e",X"d8",X"d8",X"d8",X"d8",X"d8",X"00",X"6a",X"01",X"01",X"01",
        X"01",X"00",X"00",X"b2",X"00",X"00",X"31",X"31",X"31",X"00",X"00",X"b2",X"00",X"00",X"01",X"01",
        X"00",X"00",X"5a",X"5a",X"c7",X"b2",X"d8",X"d8",X"d8",X"b2",X"9a",X"5a",X"5a",X"00",X"00",X"01",
        X"00",X"5a",X"5a",X"5a",X"5a",X"9a",X"b2",X"b2",X"b2",X"c7",X"5a",X"5a",X"5a",X"5a",X"00",X"01",
        X"00",X"5a",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"5a",X"00",X"01",
        X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"2e",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"6a",X"6a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"a5",X"01",
        X"6a",X"a5",X"21",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"2e",X"2e",X"2e",X"31",X"2e",X"2e",X"2e",X"31",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"2e",X"00",X"2e",X"31",X"2e",X"00",X"2e",X"31",X"4e",X"21",X"6a",X"01",
        X"01",X"6a",X"4e",X"31",X"2e",X"2e",X"2e",X"31",X"2e",X"2e",X"2e",X"31",X"5a",X"5a",X"5a",X"01",
        X"01",X"6a",X"4e",X"31",X"31",X"2e",X"31",X"31",X"31",X"31",X"31",X"31",X"5a",X"5a",X"5a",X"01",
        X"5a",X"5a",X"5a",X"4e",X"4e",X"4e",X"2e",X"4e",X"4e",X"4e",X"4e",X"4e",X"5a",X"5a",X"5a",X"01",
        X"5a",X"5a",X"5a",X"00",X"6a",X"6a",X"2e",X"2e",X"6a",X"6a",X"6a",X"00",X"c7",X"9a",X"6a",X"01",
        X"5a",X"5a",X"5a",X"00",X"b2",X"b2",X"2e",X"2e",X"d8",X"2e",X"d8",X"b2",X"9a",X"6a",X"01",X"01",
        X"01",X"01",X"6a",X"00",X"b2",X"d8",X"d8",X"d8",X"d8",X"d8",X"d8",X"00",X"6a",X"01",X"01",X"01",
        X"01",X"5a",X"5a",X"5a",X"00",X"00",X"31",X"31",X"31",X"00",X"00",X"b2",X"00",X"00",X"01",X"01",
        X"5a",X"5a",X"5a",X"5a",X"5a",X"b2",X"d8",X"d8",X"d8",X"b2",X"9a",X"6a",X"00",X"00",X"00",X"01",
        X"5a",X"5a",X"5a",X"5a",X"5a",X"5a",X"b2",X"b2",X"b2",X"c7",X"9a",X"5a",X"5a",X"00",X"00",X"01",
        X"00",X"5a",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"9a",X"5a",X"5a",X"5a",X"5a",X"00",X"01",
        X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"5a",X"00",X"01",
        X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"01",
        X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"2e",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"6a",X"6a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"a5",X"01",
        X"6a",X"a5",X"21",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"2e",X"2e",X"2e",X"31",X"2e",X"2e",X"2e",X"31",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"2e",X"00",X"2e",X"31",X"2e",X"00",X"2e",X"31",X"4e",X"21",X"6a",X"01",
        X"5a",X"5a",X"5a",X"31",X"2e",X"2e",X"2e",X"31",X"2e",X"2e",X"2e",X"31",X"4e",X"a5",X"01",X"01",
        X"5a",X"5a",X"5a",X"31",X"31",X"2e",X"31",X"31",X"31",X"31",X"31",X"31",X"4e",X"6a",X"01",X"01",
        X"5a",X"5a",X"5a",X"4e",X"2e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"5a",X"5a",X"5a",X"01",
        X"6a",X"c7",X"2e",X"2e",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"00",X"5a",X"5a",X"5a",X"01",
        X"01",X"6a",X"2e",X"2e",X"b2",X"b2",X"d8",X"d8",X"d8",X"2e",X"d8",X"b2",X"5a",X"5a",X"5a",X"01",
        X"01",X"01",X"6a",X"00",X"b2",X"d8",X"d8",X"d8",X"d8",X"d8",X"d8",X"00",X"6a",X"01",X"01",X"01",
        X"01",X"00",X"00",X"b2",X"00",X"00",X"31",X"31",X"31",X"00",X"00",X"5a",X"5a",X"5a",X"01",X"01",
        X"00",X"00",X"00",X"6a",X"c7",X"b2",X"d8",X"d8",X"d8",X"b2",X"5a",X"5a",X"5a",X"5a",X"5a",X"01",
        X"00",X"00",X"5a",X"5a",X"9a",X"9a",X"b2",X"b2",X"b2",X"5a",X"5a",X"5a",X"5a",X"5a",X"5a",X"01",
        X"00",X"5a",X"5a",X"5a",X"5a",X"9a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"5a",X"00",X"01",
        X"00",X"5a",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",
        X"01",X"00",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"2e",X"5a",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"5a",X"5a",X"01",
        X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"5a",X"5a",X"01",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"6a",X"6a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"a5",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"21",X"a5",X"01",
        X"01",X"4e",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"4e",X"21",X"a5",X"6a",X"01",
        X"01",X"4e",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"4e",X"21",X"6a",X"5a",X"5a",
        X"01",X"4e",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"4e",X"6a",X"5a",X"5a",X"5a",
        X"01",X"01",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"00",X"c7",X"5a",X"5a",X"5a",
        X"01",X"5a",X"5a",X"00",X"b2",X"b2",X"d8",X"d8",X"d8",X"2e",X"d8",X"b2",X"9a",X"9a",X"01",X"01",
        X"01",X"5a",X"5a",X"00",X"b2",X"d8",X"d8",X"d8",X"d8",X"d8",X"d8",X"00",X"9a",X"01",X"01",X"01",
        X"01",X"01",X"00",X"b2",X"00",X"31",X"31",X"31",X"00",X"00",X"00",X"b2",X"00",X"01",X"01",X"01",
        X"01",X"00",X"c7",X"9a",X"b2",X"b2",X"d8",X"d8",X"d8",X"d8",X"b2",X"9a",X"9a",X"00",X"01",X"01",
        X"01",X"00",X"9a",X"9a",X"9a",X"b2",X"b2",X"d8",X"d8",X"b2",X"c7",X"9a",X"9a",X"00",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"01",X"01",
        X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"21",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"6a",X"6a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"21",X"21",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"21",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"a5",X"01",
        X"6a",X"a5",X"21",X"4e",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"4e",X"a5",X"01",
        X"6a",X"a5",X"21",X"4e",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"4e",X"6a",X"01",
        X"5a",X"5a",X"5a",X"4e",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"4e",X"6a",X"01",
        X"5a",X"5a",X"5a",X"a5",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"a5",X"01",X"01",
        X"5a",X"5a",X"5a",X"6a",X"a5",X"a5",X"a5",X"a5",X"a5",X"a5",X"a5",X"a5",X"a5",X"01",X"01",X"01",
        X"6a",X"c7",X"9a",X"00",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"00",X"5a",X"5a",X"01",X"01",
        X"01",X"6a",X"9a",X"00",X"b2",X"b2",X"d8",X"d8",X"d8",X"2e",X"d8",X"b2",X"5a",X"5a",X"01",X"01",
        X"01",X"01",X"6a",X"00",X"b2",X"d8",X"d8",X"d8",X"d8",X"d8",X"d8",X"00",X"a5",X"01",X"01",X"01",
        X"01",X"01",X"01",X"b2",X"00",X"00",X"00",X"31",X"31",X"31",X"00",X"b2",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"c7",X"b2",X"b2",X"d8",X"d8",X"d8",X"d8",X"b2",X"9a",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"9a",X"9a",X"b2",X"b2",X"d8",X"d8",X"b2",X"c7",X"9a",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"9a",X"9a",X"5a",X"01",X"01",X"5a",X"9a",X"5a",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"5a",X"5a",X"5a",X"00",X"00",X"5a",X"5a",X"5a",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"00",X"2e",X"5a",X"5a",X"00",X"00",X"5a",X"5a",X"2e",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"00",X"5a",X"5a",X"00",X"00",X"00",X"00",X"5a",X"5a",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"2e",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",
        X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01",
        X"6a",X"6a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"a5",X"01",
        X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"21",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"a5",X"01",
        X"6a",X"a5",X"4e",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"4e",X"21",X"6a",X"01",
        X"01",X"6a",X"4e",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"4e",X"a5",X"01",X"01",
        X"01",X"6a",X"4e",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"4e",X"6a",X"01",X"01",
        X"01",X"01",X"6a",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"6a",X"01",X"01",X"01",
        X"01",X"6a",X"9a",X"00",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"00",X"c7",X"6a",X"01",X"01",
        X"01",X"c7",X"9a",X"00",X"b2",X"b2",X"d8",X"d8",X"d8",X"2e",X"d8",X"b2",X"9a",X"9a",X"01",X"01",
        X"01",X"5a",X"5a",X"00",X"b2",X"d8",X"d8",X"d8",X"d8",X"d8",X"d8",X"00",X"5a",X"5a",X"01",X"01",
        X"01",X"5a",X"5a",X"b2",X"00",X"00",X"31",X"31",X"31",X"00",X"00",X"b2",X"5a",X"5a",X"01",X"01",
        X"01",X"01",X"01",X"c7",X"b2",X"b2",X"d8",X"d8",X"d8",X"d8",X"b2",X"c7",X"01",X"01",X"01",X"01",
        X"01",X"01",X"00",X"9a",X"9a",X"b2",X"b2",X"d8",X"d8",X"b2",X"9a",X"9a",X"00",X"01",X"01",X"01",
        X"01",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"c7",X"9a",X"9a",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"2e",X"00",X"00",X"00",X"5a",X"5a",X"2e",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01",
        X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
        X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
        X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01", others=>X"01");
        
    constant up0 : bomberman_bitmap_type := 
       ((X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01"),
        (X"6a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01"),
        (X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"5a",X"5a",X"21",X"21",X"21",X"21",X"21",X"a5",X"01"),
        (X"6a",X"a5",X"21",X"21",X"21",X"21",X"5a",X"5a",X"2e",X"5a",X"21",X"21",X"21",X"21",X"a5",X"01"),
        (X"6a",X"a5",X"a5",X"21",X"21",X"a5",X"5a",X"5a",X"5a",X"5a",X"21",X"21",X"21",X"21",X"a5",X"01"),
        (X"6a",X"6a",X"a5",X"21",X"21",X"a5",X"a5",X"5a",X"5a",X"a5",X"21",X"21",X"21",X"a5",X"6a",X"01"),
        (X"01",X"6a",X"a5",X"a5",X"21",X"21",X"a5",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01"),
        (X"01",X"6a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01",X"01"),
        (X"01",X"01",X"6a",X"6a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"a5",X"6a",X"6a",X"01",X"01",X"01"),
        (X"01",X"6a",X"9a",X"00",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"b2",X"c7",X"6a",X"01",X"01"),
        (X"01",X"c7",X"9a",X"00",X"b2",X"b2",X"b2",X"d8",X"d8",X"2e",X"d8",X"b2",X"9a",X"9a",X"01",X"01"),
        (X"01",X"5a",X"5a",X"00",X"b2",X"b2",X"d8",X"d8",X"d8",X"d8",X"d8",X"00",X"5a",X"5a",X"01",X"01"),
        (X"01",X"5a",X"5a",X"b2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"b2",X"5a",X"5a",X"01",X"01"),
        (X"01",X"01",X"01",X"c7",X"b2",X"b2",X"b2",X"d8",X"d8",X"d8",X"b2",X"c7",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"9a",X"9a",X"b2",X"b2",X"b2",X"b2",X"b2",X"9a",X"9a",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"c7",X"9a",X"9a",X"00",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"01",X"01"),
        (X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01"),
        (X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01"),
        (X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01"),
        (X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"));
    
    constant up1 : bomberman_bitmap_type := 
       ((X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"5a",X"5a",X"a5",X"01",X"01"),
        (X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"5a",X"5a",X"2e",X"5a",X"a5",X"01"),
        (X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"5a",X"5a",X"5a",X"5a",X"a5",X"01"),
        (X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"a5",X"5a",X"5a",X"a5",X"a5",X"01"),
        (X"6a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"a5",X"a5",X"a5",X"6a",X"01"),
        (X"6a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01"),
        (X"01",X"6a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01",X"01"),
        (X"01",X"9a",X"6a",X"6a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"a5",X"a5",X"6a",X"01",X"01",X"01"),
        (X"01",X"9a",X"9a",X"00",X"00",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"c7",X"9a",X"6a",X"01",X"01"),
        (X"01",X"6a",X"9a",X"00",X"b2",X"b2",X"b2",X"d8",X"d8",X"2e",X"d8",X"9a",X"9a",X"9a",X"01",X"01"),
        (X"01",X"01",X"6a",X"00",X"b2",X"b2",X"d8",X"d8",X"d8",X"d8",X"d8",X"5a",X"2e",X"5a",X"01",X"01"),
        (X"01",X"01",X"01",X"b2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"01",X"01"),
        (X"01",X"01",X"01",X"9a",X"b2",X"b2",X"b2",X"d8",X"d8",X"d8",X"b2",X"5a",X"5a",X"5a",X"01",X"01"),
        (X"01",X"01",X"00",X"c7",X"9a",X"b2",X"b2",X"b2",X"d8",X"b2",X"c7",X"6a",X"01",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"01",X"01",X"01"),
        (X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01"),
        (X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01"),
        (X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"));
    
    constant up2 : bomberman_bitmap_type := 
       ((X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01"),
        (X"01",X"6a",X"5a",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01"),
        (X"6a",X"5a",X"5a",X"2e",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01"),
        (X"6a",X"5a",X"5a",X"5a",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01"),
        (X"6a",X"a5",X"5a",X"5a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01"),
        (X"6a",X"6a",X"a5",X"a5",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01"),
        (X"6a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01"),
        (X"01",X"6a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01",X"01"),
        (X"01",X"01",X"6a",X"6a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"a5",X"a5",X"6a",X"9a",X"01",X"01"),
        (X"01",X"6a",X"c7",X"9a",X"00",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"b2",X"c7",X"9a",X"01",X"01"),
        (X"01",X"9a",X"9a",X"9a",X"b2",X"b2",X"b2",X"d8",X"d8",X"2e",X"d8",X"b2",X"9a",X"6a",X"01",X"01"),
        (X"01",X"5a",X"2e",X"5a",X"b2",X"b2",X"d8",X"d8",X"d8",X"d8",X"d8",X"00",X"6a",X"01",X"01",X"01"),
        (X"01",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"b2",X"01",X"01",X"01",X"01"),
        (X"01",X"5a",X"5a",X"5a",X"b2",X"b2",X"b2",X"d8",X"d8",X"d8",X"b2",X"c7",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"00",X"6a",X"c7",X"b2",X"b2",X"b2",X"d8",X"b2",X"9a",X"9a",X"01",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"c7",X"9a",X"9a",X"00",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"01",X"01"),
        (X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"01",X"01"),
        (X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01"),
        (X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"));
    
    constant right0 : bomberman_bitmap_type := 
       ((X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"5a",X"5a",X"2e",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"5a",X"5a",X"5a",X"5a",X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01"),
        (X"01",X"5a",X"5a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01"),
        (X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"21",X"a5"),
        (X"01",X"01",X"6a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"4e"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"4e",X"31",X"01"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"31",X"00",X"31",X"01"),
        (X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"31",X"00",X"31",X"01"),
        (X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"31",X"00",X"31",X"4e"),
        (X"01",X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"31",X"00",X"4e",X"01"),
        (X"01",X"01",X"01",X"6a",X"a5",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"4e",X"4e",X"6a",X"01"),
        (X"01",X"01",X"01",X"01",X"b2",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"b2",X"d8",X"b2",X"c7",X"9a",X"9a",X"b2",X"2e",X"b2",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"00",X"d8",X"b2",X"9a",X"9a",X"9a",X"d8",X"d8",X"31",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"b2",X"00",X"00",X"5a",X"2e",X"5a",X"00",X"00",X"b2",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"00",X"b2",X"b2",X"5a",X"5a",X"5a",X"d8",X"b2",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"00",X"00",X"00",X"b2",X"5a",X"5a",X"5a",X"b2",X"5a",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"00",X"00",X"00",X"00",X"5a",X"c7",X"9a",X"9a",X"5a",X"5a",X"00",X"00",X"01",X"01"),
        (X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"00",X"01",X"01"),
        (X"01",X"01",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"2e",X"5a",X"00",X"00",X"01",X"01"),
        (X"01",X"01",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01"),
        (X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"));
    
    constant right1 : bomberman_bitmap_type := 
       ((X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"5a",X"5a",X"2e",X"5a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01"),
        (X"5a",X"5a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"4e",X"01"),
        (X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"4e",X"4e",X"01",X"01"),
        (X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"4e",X"4e",X"4e",X"31",X"00",X"01",X"01"),
        (X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"4e",X"31",X"31",X"00",X"31",X"31",X"00",X"01",X"01"),
        (X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"4e",X"31",X"31",X"00",X"31",X"31",X"00",X"01",X"01"),
        (X"01",X"a5",X"a5",X"21",X"21",X"21",X"21",X"4e",X"31",X"31",X"00",X"31",X"31",X"00",X"4e",X"01"),
        (X"01",X"6a",X"a5",X"a5",X"a5",X"21",X"21",X"4e",X"31",X"31",X"00",X"31",X"4e",X"4e",X"01",X"01"),
        (X"01",X"01",X"6a",X"6a",X"a5",X"a5",X"a5",X"6a",X"4e",X"4e",X"4e",X"4e",X"6a",X"6a",X"01",X"01"),
        (X"01",X"01",X"5a",X"00",X"00",X"6a",X"6a",X"6a",X"6a",X"6a",X"5a",X"2e",X"5a",X"01",X"01",X"01"),
        (X"01",X"01",X"5a",X"b2",X"b2",X"d8",X"b2",X"c7",X"9a",X"9a",X"5a",X"5a",X"5a",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"00",X"b2",X"d8",X"b2",X"b2",X"9a",X"9a",X"5a",X"5a",X"5a",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"b2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"b2",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"00",X"b2",X"b2",X"9a",X"9a",X"d8",X"b2",X"b2",X"c7",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"00",X"00",X"5a",X"c7",X"9a",X"9a",X"6a",X"b2",X"6a",X"9a",X"9a",X"5a",X"5a",X"01"),
        (X"01",X"00",X"00",X"5a",X"5a",X"9a",X"9a",X"6a",X"00",X"00",X"6a",X"6a",X"5a",X"5a",X"5a",X"01"),
        (X"01",X"00",X"00",X"5a",X"5a",X"5a",X"6a",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"01"),
        (X"01",X"00",X"00",X"5a",X"5a",X"2e",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"00",X"00",X"00"),
        (X"01",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01"),
        (X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01"),
        (X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"));
    
    constant right2 : bomberman_bitmap_type := 
       ((X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01"),
        (X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01"),
        (X"01",X"5a",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"4e"),
        (X"5a",X"5a",X"2e",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e"),
        (X"5a",X"5a",X"5a",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e"),
        (X"01",X"5a",X"5a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"4e"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"01"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"4e",X"01"),
        (X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"4e",X"01"),
        (X"01",X"01",X"01",X"6a",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"a5",X"6a",X"5a",X"5a"),
        (X"01",X"01",X"01",X"01",X"00",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"b2",X"6a",X"5a",X"5a"),
        (X"01",X"01",X"01",X"01",X"b2",X"00",X"b2",X"9a",X"9a",X"b2",X"2e",X"d8",X"b2",X"6a",X"5a",X"5a"),
        (X"01",X"01",X"01",X"01",X"b2",X"b2",X"c7",X"9a",X"b2",X"d8",X"d8",X"b2",X"31",X"01",X"01",X"01"),
        (X"01",X"01",X"00",X"6a",X"5a",X"2e",X"5a",X"9a",X"00",X"00",X"00",X"00",X"b2",X"00",X"01",X"01"),
        (X"01",X"00",X"6a",X"c7",X"5a",X"5a",X"5a",X"6a",X"b2",X"9a",X"c7",X"b2",X"00",X"00",X"00",X"01"),
        (X"00",X"00",X"5a",X"9a",X"5a",X"5a",X"5a",X"b2",X"6a",X"9a",X"9a",X"9a",X"6a",X"5a",X"5a",X"00"),
        (X"00",X"00",X"5a",X"5a",X"9a",X"00",X"00",X"00",X"00",X"6a",X"9a",X"9a",X"5a",X"2e",X"5a",X"00"),
        (X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"9a",X"5a",X"5a",X"5a",X"00",X"00"),
        (X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00"),
        (X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"00",X"00",X"00",X"01"),
        (X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"));
    
    constant down0 : bomberman_bitmap_type := 
       ((X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"2e",X"5a",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01"),
        (X"6a",X"6a",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"a5",X"01"),
        (X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01"),
        (X"6a",X"a5",X"21",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"a5",X"01"),
        (X"6a",X"a5",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"a5",X"01"),
        (X"6a",X"a5",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"6a",X"01"),
        (X"01",X"6a",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"a5",X"01",X"01"),
        (X"01",X"6a",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"6a",X"01",X"01"),
        (X"01",X"01",X"6a",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"6a",X"01",X"01",X"01"),
        (X"01",X"6a",X"9a",X"00",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"00",X"c7",X"6a",X"01",X"01"),
        (X"01",X"c7",X"9a",X"00",X"b2",X"b2",X"d8",X"d8",X"d8",X"2e",X"d8",X"b2",X"9a",X"9a",X"01",X"01"),
        (X"01",X"5a",X"5a",X"00",X"b2",X"d8",X"d8",X"d8",X"d8",X"d8",X"d8",X"00",X"5a",X"5a",X"01",X"01"),
        (X"01",X"5a",X"5a",X"b2",X"00",X"00",X"31",X"31",X"31",X"00",X"00",X"b2",X"5a",X"5a",X"01",X"01"),
        (X"01",X"01",X"01",X"c7",X"b2",X"b2",X"d8",X"d8",X"d8",X"d8",X"b2",X"c7",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"00",X"9a",X"9a",X"b2",X"b2",X"d8",X"d8",X"b2",X"9a",X"9a",X"00",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"c7",X"9a",X"9a",X"00",X"00",X"01",X"01"),
        (X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01"),
        (X"01",X"00",X"00",X"5a",X"5a",X"2e",X"00",X"00",X"00",X"5a",X"5a",X"2e",X"00",X"00",X"01",X"01"),
        (X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01"),
        (X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01"),
        (X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"));
    
    constant down1 : bomberman_bitmap_type := 
       ((X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"5a",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"5a",X"5a",X"2e",X"5a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"5a",X"5a",X"5a",X"5a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"5a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01"),
        (X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01"),
        (X"6a",X"a5",X"21",X"21",X"21",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"21",X"a5",X"01"),
        (X"6a",X"a5",X"a5",X"21",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"4e",X"a5",X"01"),
        (X"6a",X"a5",X"a5",X"21",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"4e",X"a5",X"01"),
        (X"6a",X"6a",X"a5",X"a5",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"4e",X"6a",X"01"),
        (X"01",X"6a",X"6a",X"a5",X"4e",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"4e",X"6a",X"01"),
        (X"01",X"01",X"6a",X"6a",X"6a",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"6a",X"01",X"01"),
        (X"01",X"6a",X"9a",X"00",X"00",X"6a",X"6a",X"6a",X"6a",X"5a",X"2e",X"5a",X"c7",X"9a",X"01",X"01"),
        (X"01",X"9a",X"9a",X"00",X"b2",X"b2",X"d8",X"d8",X"b2",X"5a",X"5a",X"5a",X"9a",X"6a",X"01",X"01"),
        (X"01",X"5a",X"5a",X"00",X"b2",X"d8",X"d8",X"d8",X"b2",X"5a",X"5a",X"5a",X"6a",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"9a",X"00",X"00",X"31",X"31",X"31",X"00",X"00",X"6a",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"00",X"c7",X"9a",X"b2",X"d8",X"d8",X"d8",X"b2",X"9a",X"6a",X"00",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"9a",X"9a",X"9a",X"b2",X"d8",X"b2",X"c7",X"9a",X"5a",X"00",X"00",X"01",X"01"),
        (X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01"),
        (X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"5a",X"00",X"00",X"01",X"01",X"01"),
        (X"00",X"00",X"5a",X"5a",X"2e",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01"),
        (X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"));
    
    constant down2 : bomberman_bitmap_type := 
       ((X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"2e",X"5a",X"01"),
        (X"01",X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"a5",X"5a",X"5a",X"5a",X"5a",X"01"),
        (X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"5a",X"01",X"01"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01"),
        (X"01",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"01",X"01"),
        (X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01"),
        (X"6a",X"a5",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"21",X"21",X"a5",X"01"),
        (X"6a",X"4e",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"21",X"21",X"a5",X"01"),
        (X"6a",X"4e",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"21",X"21",X"a5",X"01"),
        (X"6a",X"4e",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"21",X"a5",X"6a",X"01"),
        (X"6a",X"4e",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"a5",X"6a",X"01",X"01"),
        (X"01",X"6a",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"4e",X"6a",X"6a",X"6a",X"01",X"01",X"01"),
        (X"01",X"9a",X"9a",X"5a",X"2e",X"5a",X"6a",X"6a",X"6a",X"6a",X"b2",X"b2",X"c7",X"6a",X"01",X"01"),
        (X"01",X"6a",X"9a",X"5a",X"5a",X"5a",X"b2",X"b2",X"d8",X"2e",X"d8",X"b2",X"9a",X"9a",X"01",X"01"),
        (X"01",X"01",X"6a",X"5a",X"5a",X"5a",X"b2",X"b2",X"d8",X"d8",X"d8",X"00",X"5a",X"5a",X"01",X"01"),
        (X"01",X"01",X"01",X"6a",X"00",X"00",X"31",X"31",X"31",X"00",X"00",X"c7",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"00",X"6a",X"c7",X"b2",X"b2",X"d8",X"d8",X"b2",X"9a",X"9a",X"01",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"5a",X"9a",X"9a",X"b2",X"b2",X"b2",X"c7",X"9a",X"9a",X"00",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"01",X"01"),
        (X"01",X"00",X"00",X"00",X"5a",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01",X"01"),
        (X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"2e",X"5a",X"00",X"01",X"01"),
        (X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"));
    
    constant left0 : bomberman_bitmap_type := 
       ((X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"2e",X"5a"),
        (X"01",X"01",X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"01",X"5a",X"5a",X"5a",X"5a"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"5a",X"5a",X"01"),
        (X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01"),
        (X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01"),
        (X"4e",X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01"),
        (X"01",X"31",X"4e",X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01"),
        (X"01",X"31",X"00",X"31",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01"),
        (X"01",X"31",X"00",X"31",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01"),
        (X"4e",X"31",X"00",X"31",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01"),
        (X"01",X"4e",X"00",X"31",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01",X"01"),
        (X"01",X"6a",X"4e",X"4e",X"a5",X"a5",X"21",X"21",X"21",X"21",X"a5",X"6a",X"6a",X"01",X"01",X"01"),
        (X"01",X"01",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"b2",X"b2",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"b2",X"d8",X"b2",X"c7",X"9a",X"9a",X"b2",X"2e",X"d8",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"31",X"d8",X"b2",X"9a",X"9a",X"9a",X"d8",X"d8",X"00",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"b2",X"00",X"00",X"5a",X"2e",X"5a",X"00",X"00",X"b2",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"00",X"b2",X"b2",X"5a",X"5a",X"5a",X"d8",X"b2",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"00",X"00",X"5a",X"b2",X"5a",X"5a",X"5a",X"b2",X"00",X"00",X"01",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"00",X"5a",X"5a",X"c7",X"9a",X"9a",X"5a",X"00",X"00",X"00",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"00",X"00",X"00",X"9a",X"9a",X"9a",X"00",X"00",X"00",X"00",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"2e",X"5a",X"00",X"00",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"));
    
    constant left1 : bomberman_bitmap_type := 
       ((X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"a5",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01",X"01"),
        (X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01",X"01"),
        (X"4e",X"a5",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"5a",X"5a",X"01"),
        (X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"5a",X"5a",X"2e",X"5a"),
        (X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"5a",X"5a",X"5a",X"5a"),
        (X"4e",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"5a",X"5a",X"01"),
        (X"01",X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01"),
        (X"01",X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01",X"01"),
        (X"01",X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01",X"01"),
        (X"5a",X"5a",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"a5",X"6a",X"01",X"01",X"01"),
        (X"5a",X"5a",X"6a",X"b2",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"6a",X"b2",X"01",X"01",X"01",X"01"),
        (X"5a",X"5a",X"6a",X"b2",X"d8",X"b2",X"6a",X"c7",X"9a",X"b2",X"b2",X"d8",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"31",X"d8",X"b2",X"b2",X"6a",X"9a",X"9a",X"d8",X"d8",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"00",X"b2",X"00",X"00",X"00",X"00",X"9a",X"5a",X"2e",X"5a",X"6a",X"01",X"01",X"01"),
        (X"01",X"00",X"00",X"00",X"b2",X"9a",X"9a",X"b2",X"6a",X"5a",X"5a",X"5a",X"9a",X"6a",X"01",X"01"),
        (X"00",X"5a",X"5a",X"6a",X"c7",X"9a",X"9a",X"b2",X"b2",X"5a",X"5a",X"5a",X"9a",X"5a",X"00",X"01"),
        (X"00",X"5a",X"2e",X"5a",X"9a",X"9a",X"6a",X"00",X"00",X"00",X"00",X"9a",X"5a",X"5a",X"00",X"01"),
        (X"00",X"00",X"5a",X"5a",X"5a",X"9a",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"01"),
        (X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01"),
        (X"01",X"00",X"00",X"00",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01"),
        (X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"));
    
    constant left2 : bomberman_bitmap_type := 
       ((X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5a",X"5a",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"6a",X"a5",X"a5",X"21",X"21",X"21",X"a5",X"5a",X"5a",X"2e",X"5a"),
        (X"01",X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"5a",X"5a"),
        (X"01",X"01",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"2e",X"21",X"21",X"a5",X"01"),
        (X"01",X"4e",X"6a",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5",X"01"),
        (X"01",X"01",X"4e",X"4e",X"a5",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5"),
        (X"01",X"01",X"00",X"31",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"a5"),
        (X"01",X"01",X"00",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"21",X"21",X"21",X"21",X"21",X"a5"),
        (X"01",X"01",X"00",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"21",X"21",X"21",X"21",X"a5",X"6a"),
        (X"01",X"4e",X"00",X"31",X"31",X"00",X"31",X"31",X"4e",X"21",X"21",X"21",X"21",X"21",X"a5",X"01"),
        (X"01",X"6a",X"4e",X"4e",X"31",X"00",X"31",X"31",X"4e",X"21",X"21",X"21",X"21",X"a5",X"6a",X"01"),
        (X"01",X"01",X"6a",X"6a",X"4e",X"4e",X"4e",X"4e",X"21",X"21",X"21",X"a5",X"6a",X"6a",X"01",X"01"),
        (X"01",X"01",X"01",X"5a",X"2e",X"5a",X"6a",X"6a",X"6a",X"6a",X"6a",X"b2",X"b2",X"5a",X"01",X"01"),
        (X"01",X"01",X"01",X"5a",X"5a",X"5a",X"c7",X"9a",X"9a",X"b2",X"d8",X"2e",X"d8",X"5a",X"01",X"01"),
        (X"01",X"01",X"01",X"5a",X"5a",X"5a",X"9a",X"9a",X"b2",X"b2",X"d8",X"d8",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"b2",X"31",X"00",X"00",X"00",X"00",X"00",X"00",X"b2",X"01",X"01",X"01"),
        (X"01",X"01",X"00",X"00",X"9a",X"b2",X"b2",X"b2",X"d8",X"c7",X"9a",X"b2",X"00",X"01",X"01",X"01"),
        (X"01",X"5a",X"5a",X"c7",X"9a",X"6a",X"b2",X"b2",X"6a",X"9a",X"9a",X"9a",X"5a",X"00",X"01",X"01"),
        (X"01",X"5a",X"5a",X"5a",X"6a",X"6a",X"00",X"00",X"00",X"6a",X"9a",X"9a",X"5a",X"5a",X"00",X"01"),
        (X"01",X"00",X"5a",X"5a",X"5a",X"00",X"00",X"00",X"00",X"00",X"6a",X"5a",X"5a",X"2e",X"00",X"01"),
        (X"00",X"00",X"00",X"5a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"00",X"01"),
        (X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5a",X"5a",X"5a",X"5a",X"00",X"01"),
        (X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"));
        
   type walking_bomberman_type is array(0 to 2) of bomberman_bitmap_type;
   constant up_frames    : walking_bomberman_type := (up0, up1, up2);
   constant down_frames  : walking_bomberman_type := (down0, down1, down2);
   constant right_frames : walking_bomberman_type := (right0, right1, right2);
   constant left_frames  : walking_bomberman_type := (left0, left1, left2);
end package;