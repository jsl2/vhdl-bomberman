use work.graphics_pkg.all;

package explosions_pkg is
    -- quite inefficient blockram : 35 tiles used, but 64 available
    type explosions_rom_type is array(0 to (2**14 - 1)) of pixel_type;
    constant MAX_EXPLOSIONS : integer := 32; 
    
    constant EXPLOSION_FRAMES : explosions_rom_type := 
   (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"01",X"65",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"65",X"d7",X"d7",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"65",X"d7",X"d7",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"d7",X"99",X"99",X"d7",X"65",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"65",X"d7",X"99",X"99",X"d7",X"65",X"bd",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"bd",X"65",X"d7",X"99",X"8a",X"d7",X"65",X"bd",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"bd",X"65",X"99",X"99",X"8a",X"99",X"d7",X"bd",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"65",X"d7",X"99",X"99",X"8a",X"99",X"d7",X"65",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"d7",X"d7",X"99",X"8a",X"8a",X"8a",X"d7",X"65",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"8a",X"d7",X"65",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"65",X"65",X"d7",X"99",X"8a",X"8a",X"99",X"99",X"d7",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"d7",X"d7",X"99",X"99",X"8a",X"99",X"d7",X"d7",X"65",X"01",X"01",X"01",
    X"01",X"01",X"01",X"b4",X"65",X"d7",X"99",X"8a",X"8a",X"8a",X"99",X"d7",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"65",X"d7",X"8a",X"8a",X"2e",X"8a",X"99",X"d7",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"01",X"65",X"65",X"65",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"d7",X"d7",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"65",X"d7",X"99",X"99",X"d7",X"65",X"bd",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"65",X"d7",X"99",X"99",X"d7",X"65",X"bd",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"bd",X"d7",X"99",X"99",X"8a",X"99",X"d7",X"65",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"65",X"d7",X"99",X"8a",X"8a",X"99",X"d7",X"65",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"65",X"d7",X"99",X"8a",X"8a",X"8a",X"d7",X"65",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"65",X"99",X"99",X"8a",X"2e",X"8a",X"99",X"d7",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"65",X"d7",X"99",X"99",X"8a",X"2e",X"8a",X"99",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"8a",X"8a",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"8a",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"65",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"d7",X"d7",X"99",X"99",X"8a",X"2e",X"8a",X"99",X"d7",X"d7",X"65",X"01",X"01",
    X"01",X"01",X"b4",X"65",X"d7",X"99",X"8a",X"2e",X"8a",X"8a",X"8a",X"99",X"d7",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"65",X"d7",X"8a",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"bd",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"01",X"01",X"65",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"bd",X"01",X"65",X"bd",X"bd",X"65",X"65",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"bd",X"65",X"d7",X"65",X"65",X"d7",X"65",X"bd",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"65",X"d7",X"99",X"d7",X"d7",X"99",X"d7",X"65",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"65",X"d7",X"99",X"99",X"d7",X"99",X"d7",X"65",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"d7",X"99",X"99",X"8a",X"99",X"8a",X"99",X"d7",X"65",X"01",X"01",X"01",
    X"01",X"01",X"01",X"65",X"d7",X"99",X"8a",X"2e",X"8a",X"8a",X"99",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"8a",X"8a",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"65",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"bd",X"01",X"01",
    X"01",X"01",X"65",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"65",X"bd",X"01",
    X"01",X"bd",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"d7",X"65",X"bd",X"01",
    X"01",X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"d7",X"65",X"bd",X"01",
    X"01",X"65",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"bd",X"01",
    X"01",X"bd",X"d7",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",X"65",X"01",
    X"01",X"b4",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"99",X"d7",X"bd",X"01",
    X"01",X"bd",X"65",X"d7",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"bd",X"01",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"01",X"bd",X"01",X"01",X"65",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"01",X"65",X"bd",X"bd",X"65",X"bd",X"65",X"65",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"65",X"d7",X"65",X"d7",X"d7",X"65",X"d7",X"65",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"65",X"d7",X"99",X"d7",X"99",X"d7",X"d7",X"99",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"01",X"65",X"d7",X"99",X"99",X"8a",X"99",X"d7",X"99",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"d7",X"99",X"99",X"8a",X"8a",X"8a",X"99",X"8a",X"99",X"d7",X"65",X"01",X"01",
    X"01",X"01",X"65",X"d7",X"99",X"8a",X"2e",X"8a",X"8a",X"8a",X"8a",X"99",X"d7",X"65",X"bd",X"01",
    X"01",X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"8a",X"2e",X"8a",X"8a",X"d7",X"65",X"bd",X"01",
    X"01",X"bd",X"65",X"99",X"99",X"8a",X"2e",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"bd",X"01",
    X"01",X"65",X"d7",X"99",X"99",X"8a",X"2e",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"65",X"bd",
    X"bd",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"d7",X"65",X"bd",
    X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"d7",X"65",X"bd",
    X"65",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"bd",
    X"bd",X"d7",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",X"65",
    X"b4",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"99",X"d7",X"bd",
    X"bd",X"65",X"d7",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"bd",
    X"01",X"01",X"01",X"bd",X"65",X"01",X"bd",X"65",X"65",X"bd",X"01",X"bd",X"01",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"65",X"d7",X"65",X"65",X"d7",X"d7",X"bd",X"bd",X"65",X"bd",X"65",X"01",X"01",
    X"01",X"b4",X"65",X"65",X"d7",X"d7",X"d7",X"99",X"99",X"d7",X"65",X"d7",X"65",X"65",X"b4",X"01",
    X"01",X"bd",X"65",X"d7",X"d7",X"99",X"d7",X"99",X"8a",X"99",X"d7",X"d7",X"d7",X"65",X"bd",X"01",
    X"01",X"65",X"d7",X"d7",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"99",X"99",X"d7",X"d7",X"65",X"01",
    X"bd",X"65",X"d7",X"d7",X"99",X"8a",X"99",X"8a",X"2e",X"8a",X"8a",X"99",X"99",X"d7",X"65",X"bd",
    X"65",X"65",X"d7",X"99",X"99",X"8a",X"8a",X"2e",X"2e",X"8a",X"2e",X"8a",X"99",X"d7",X"d7",X"65",
    X"65",X"d7",X"d7",X"99",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"65",
    X"65",X"d7",X"99",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",X"65",
    X"65",X"d7",X"99",X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",
    X"d7",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",
    X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"d7",X"d7",
    X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",
    X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",
    X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"99",X"d7",
    X"65",X"d7",X"8a",X"8a",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",
    X"01",X"01",X"01",X"bd",X"65",X"d7",X"8a",X"8a",X"2e",X"8a",X"99",X"d7",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"b4",X"65",X"d7",X"99",X"8a",X"8a",X"8a",X"99",X"d7",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"d7",X"d7",X"99",X"99",X"8a",X"99",X"d7",X"d7",X"65",X"01",X"01",X"01",
    X"01",X"01",X"01",X"65",X"65",X"d7",X"99",X"8a",X"8a",X"99",X"99",X"d7",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"8a",X"d7",X"65",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"d7",X"d7",X"99",X"8a",X"8a",X"8a",X"d7",X"65",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"65",X"d7",X"99",X"99",X"8a",X"99",X"d7",X"65",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"bd",X"65",X"99",X"99",X"8a",X"99",X"d7",X"bd",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"bd",X"65",X"d7",X"99",X"8a",X"d7",X"65",X"bd",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"65",X"d7",X"99",X"99",X"d7",X"65",X"bd",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"d7",X"99",X"99",X"d7",X"65",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"65",X"d7",X"d7",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"65",X"d7",X"d7",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"01",X"65",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"bd",X"65",X"d7",X"8a",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"bd",X"01",X"01",
    X"01",X"01",X"b4",X"65",X"d7",X"99",X"8a",X"2e",X"8a",X"8a",X"8a",X"99",X"d7",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"d7",X"d7",X"99",X"99",X"8a",X"2e",X"8a",X"99",X"d7",X"d7",X"65",X"01",X"01",
    X"01",X"01",X"65",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"8a",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"8a",X"8a",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"01",X"65",X"d7",X"99",X"99",X"8a",X"2e",X"8a",X"99",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"65",X"99",X"99",X"8a",X"2e",X"8a",X"99",X"d7",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"65",X"d7",X"99",X"8a",X"8a",X"8a",X"d7",X"65",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"65",X"d7",X"99",X"8a",X"8a",X"99",X"d7",X"65",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"bd",X"d7",X"99",X"99",X"8a",X"99",X"d7",X"65",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"65",X"d7",X"99",X"99",X"d7",X"65",X"bd",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"65",X"d7",X"99",X"99",X"d7",X"65",X"bd",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"d7",X"d7",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"01",X"65",X"65",X"65",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"bd",X"65",X"d7",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"bd",X"01",
    X"01",X"b4",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"99",X"d7",X"bd",X"01",
    X"01",X"bd",X"d7",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",X"65",X"01",
    X"01",X"65",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"bd",X"01",
    X"01",X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"d7",X"65",X"bd",X"01",
    X"01",X"bd",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"d7",X"65",X"bd",X"01",
    X"01",X"01",X"65",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"65",X"bd",X"01",
    X"01",X"01",X"bd",X"65",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"8a",X"8a",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"01",X"65",X"d7",X"99",X"8a",X"2e",X"8a",X"8a",X"99",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"d7",X"99",X"99",X"8a",X"99",X"8a",X"99",X"d7",X"65",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"65",X"d7",X"99",X"99",X"d7",X"99",X"d7",X"65",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"65",X"d7",X"99",X"d7",X"d7",X"99",X"d7",X"65",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"bd",X"65",X"d7",X"65",X"65",X"d7",X"65",X"bd",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"bd",X"01",X"65",X"bd",X"bd",X"65",X"65",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"01",X"01",X"65",X"01",X"01",X"01",X"01",X"01",X"01",
    X"bd",X"65",X"d7",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"bd",
    X"b4",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"99",X"d7",X"bd",
    X"bd",X"d7",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",X"65",
    X"65",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"bd",
    X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"d7",X"65",X"bd",
    X"bd",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"d7",X"65",X"bd",
    X"01",X"65",X"d7",X"99",X"99",X"8a",X"2e",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"65",X"bd",
    X"01",X"bd",X"65",X"99",X"99",X"8a",X"2e",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"bd",X"01",
    X"01",X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"8a",X"2e",X"8a",X"8a",X"d7",X"65",X"bd",X"01",
    X"01",X"01",X"65",X"d7",X"99",X"8a",X"2e",X"8a",X"8a",X"8a",X"8a",X"99",X"d7",X"65",X"bd",X"01",
    X"01",X"01",X"bd",X"d7",X"99",X"99",X"8a",X"8a",X"8a",X"99",X"8a",X"99",X"d7",X"65",X"01",X"01",
    X"01",X"01",X"01",X"65",X"d7",X"99",X"99",X"8a",X"99",X"d7",X"99",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"01",X"65",X"d7",X"99",X"d7",X"99",X"d7",X"d7",X"99",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"65",X"d7",X"65",X"d7",X"d7",X"65",X"d7",X"65",X"bd",X"01",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"01",X"65",X"bd",X"bd",X"65",X"bd",X"65",X"65",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"01",X"bd",X"01",X"01",X"65",X"01",X"01",X"01",X"01",X"01",
    X"65",X"d7",X"8a",X"8a",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",
    X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"99",X"d7",
    X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",
    X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",
    X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"d7",X"d7",
    X"d7",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",
    X"65",X"d7",X"99",X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",
    X"65",X"d7",X"99",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",X"65",
    X"65",X"d7",X"d7",X"99",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"65",
    X"65",X"65",X"d7",X"99",X"99",X"8a",X"8a",X"2e",X"2e",X"8a",X"2e",X"8a",X"99",X"d7",X"d7",X"65",
    X"bd",X"65",X"d7",X"d7",X"99",X"8a",X"99",X"8a",X"2e",X"8a",X"8a",X"99",X"99",X"d7",X"65",X"bd",
    X"01",X"65",X"d7",X"d7",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"99",X"99",X"d7",X"d7",X"65",X"01",
    X"01",X"bd",X"65",X"d7",X"d7",X"99",X"d7",X"99",X"8a",X"99",X"d7",X"d7",X"d7",X"65",X"bd",X"01",
    X"01",X"b4",X"65",X"65",X"d7",X"d7",X"d7",X"99",X"99",X"d7",X"65",X"d7",X"65",X"65",X"b4",X"01",
    X"01",X"01",X"bd",X"65",X"d7",X"65",X"65",X"d7",X"d7",X"bd",X"bd",X"65",X"bd",X"65",X"01",X"01",
    X"01",X"01",X"01",X"bd",X"65",X"01",X"bd",X"65",X"65",X"bd",X"01",X"bd",X"01",X"bd",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"bd",X"b4",X"b4",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"bd",X"bd",X"65",X"b4",X"b4",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"65",X"65",X"d7",X"65",X"65",X"d7",X"65",X"65",
    X"01",X"01",X"b4",X"bd",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",
    X"01",X"bd",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"8a",
    X"bd",X"65",X"65",X"d7",X"d7",X"99",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",
    X"01",X"bd",X"65",X"d7",X"d7",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"2e",X"8a",X"8a",X"8a",X"2e",
    X"bd",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"99",X"99",X"99",X"99",X"8a",X"99",X"99",X"8a",X"8a",
    X"01",X"01",X"b4",X"bd",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"99",X"d7",X"99",X"d7",X"99",X"99",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"65",X"d7",X"65",X"65",X"65",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"bd",X"bd",X"b4",X"b4",X"bd",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"bd",X"bd",X"b4",X"b4",X"bd",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"65",X"d7",X"65",X"65",X"65",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",
    X"01",X"01",X"b4",X"bd",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"99",X"d7",X"99",X"d7",X"99",X"99",
    X"bd",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"99",X"99",X"99",X"99",X"8a",X"99",X"99",X"8a",X"8a",
    X"01",X"bd",X"65",X"d7",X"d7",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"2e",X"8a",X"8a",X"8a",X"2e",
    X"bd",X"65",X"d7",X"d7",X"99",X"8a",X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",
    X"65",X"d7",X"d7",X"d7",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"8a",X"8a",X"2e",X"2e",X"8a",X"2e",
    X"bd",X"65",X"65",X"d7",X"d7",X"99",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",
    X"01",X"bd",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"8a",
    X"01",X"01",X"b4",X"bd",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"65",X"65",X"d7",X"65",X"65",X"d7",X"65",X"65",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"bd",X"bd",X"65",X"b4",X"b4",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"bd",X"b4",X"b4",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"bd",X"b4",X"b4",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"bd",X"bd",X"65",X"b4",X"b4",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"65",X"65",X"d7",X"65",X"65",X"d7",X"65",X"65",
    X"01",X"01",X"b4",X"bd",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",
    X"01",X"bd",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"8a",
    X"bd",X"65",X"65",X"d7",X"d7",X"99",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",
    X"65",X"d7",X"d7",X"d7",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"8a",X"8a",X"2e",X"2e",X"8a",X"2e",
    X"01",X"65",X"d7",X"99",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",
    X"01",X"bd",X"65",X"d7",X"99",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"bd",X"65",X"d7",X"d7",X"99",X"8a",X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",
    X"01",X"bd",X"65",X"d7",X"d7",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"2e",X"8a",X"8a",X"8a",X"2e",
    X"bd",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"99",X"99",X"99",X"99",X"8a",X"99",X"99",X"8a",X"8a",
    X"01",X"01",X"b4",X"bd",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"99",X"d7",X"99",X"d7",X"99",X"99",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"65",X"d7",X"65",X"65",X"65",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"bd",X"bd",X"b4",X"b4",X"bd",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"65",X"d7",X"65",X"65",X"65",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",
    X"01",X"01",X"b4",X"bd",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"99",X"d7",X"99",X"d7",X"99",X"99",
    X"bd",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"99",X"99",X"99",X"99",X"8a",X"99",X"99",X"8a",X"8a",
    X"01",X"bd",X"65",X"d7",X"d7",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"2e",X"8a",X"8a",X"8a",X"2e",
    X"bd",X"65",X"d7",X"d7",X"99",X"99",X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",
    X"01",X"bd",X"65",X"d7",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"bd",X"bd",X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"bd",X"65",X"d7",X"99",X"99",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"01",X"65",X"d7",X"99",X"99",X"8a",X"8a",X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",
    X"65",X"d7",X"d7",X"d7",X"99",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"8a",X"2e",X"2e",X"8a",X"2e",
    X"bd",X"65",X"65",X"d7",X"d7",X"d7",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",
    X"01",X"bd",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"8a",
    X"01",X"01",X"b4",X"bd",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"65",X"65",X"d7",X"65",X"65",X"d7",X"65",X"65",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"bd",X"bd",X"65",X"b4",X"b4",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"65",X"65",X"d7",X"65",X"65",X"d7",X"65",X"65",
    X"01",X"01",X"b4",X"bd",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",
    X"01",X"bd",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"8a",
    X"bd",X"65",X"65",X"d7",X"d7",X"d7",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",
    X"65",X"d7",X"d7",X"d7",X"99",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"8a",X"2e",X"2e",X"8a",X"2e",
    X"01",X"65",X"d7",X"99",X"99",X"8a",X"8a",X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",
    X"bd",X"65",X"d7",X"d7",X"99",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"65",X"d7",X"99",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"bd",X"bd",X"d7",X"99",X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"01",X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"bd",X"65",X"d7",X"d7",X"99",X"99",X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",
    X"01",X"bd",X"65",X"d7",X"d7",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"2e",X"8a",X"8a",X"8a",X"2e",
    X"bd",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"99",X"99",X"99",X"99",X"8a",X"99",X"99",X"8a",X"8a",
    X"01",X"01",X"b4",X"bd",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"99",X"d7",X"99",X"d7",X"99",X"99",
    X"01",X"01",X"01",X"01",X"01",X"bd",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"b4",X"b4",X"bd",X"bd",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"b4",X"b4",X"65",X"bd",X"bd",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"65",X"65",X"d7",X"65",X"65",X"d7",X"65",X"65",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",
    X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"65",X"bd",X"b4",X"01",X"01",
    X"8a",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"bd",X"01",
    X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"99",X"99",X"99",X"99",X"d7",X"d7",X"65",X"65",X"bd",
    X"2e",X"8a",X"8a",X"8a",X"2e",X"8a",X"8a",X"8a",X"99",X"99",X"99",X"d7",X"d7",X"65",X"bd",X"01",
    X"8a",X"8a",X"99",X"99",X"8a",X"99",X"99",X"99",X"99",X"d7",X"d7",X"d7",X"65",X"65",X"65",X"bd",
    X"99",X"99",X"d7",X"99",X"d7",X"99",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"bd",X"b4",X"01",X"01",
    X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",
    X"65",X"65",X"65",X"d7",X"65",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"bd",X"b4",X"b4",X"bd",X"bd",X"bd",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"bd",X"b4",X"b4",X"bd",X"bd",X"bd",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"65",X"65",X"65",X"d7",X"65",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",
    X"99",X"99",X"d7",X"99",X"d7",X"99",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"bd",X"b4",X"01",X"01",
    X"8a",X"8a",X"99",X"99",X"8a",X"99",X"99",X"99",X"99",X"d7",X"d7",X"d7",X"65",X"65",X"65",X"bd",
    X"2e",X"8a",X"8a",X"8a",X"2e",X"8a",X"8a",X"8a",X"99",X"99",X"99",X"d7",X"d7",X"65",X"bd",X"01",
    X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"8a",X"99",X"d7",X"d7",X"65",X"bd",
    X"2e",X"8a",X"2e",X"2e",X"8a",X"8a",X"8a",X"8a",X"8a",X"99",X"99",X"99",X"d7",X"d7",X"d7",X"65",
    X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"99",X"99",X"99",X"99",X"d7",X"d7",X"65",X"65",X"bd",
    X"8a",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"bd",X"01",
    X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"65",X"bd",X"b4",X"01",X"01",
    X"65",X"65",X"d7",X"65",X"65",X"d7",X"65",X"65",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",
    X"b4",X"b4",X"65",X"bd",X"bd",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"b4",X"b4",X"bd",X"bd",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"b4",X"b4",X"bd",X"bd",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"b4",X"b4",X"65",X"bd",X"bd",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"65",X"65",X"d7",X"65",X"65",X"d7",X"65",X"65",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",
    X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"65",X"bd",X"b4",X"01",X"01",
    X"8a",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"bd",X"01",
    X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"99",X"99",X"99",X"99",X"d7",X"d7",X"65",X"65",X"bd",
    X"2e",X"8a",X"2e",X"2e",X"8a",X"8a",X"8a",X"8a",X"8a",X"99",X"99",X"99",X"d7",X"d7",X"d7",X"65",
    X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"99",X"d7",X"65",X"01",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"99",X"d7",X"65",X"bd",X"01",
    X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"8a",X"99",X"d7",X"d7",X"65",X"bd",
    X"2e",X"8a",X"8a",X"8a",X"2e",X"8a",X"8a",X"8a",X"99",X"99",X"99",X"d7",X"d7",X"65",X"bd",X"01",
    X"8a",X"8a",X"99",X"99",X"8a",X"99",X"99",X"99",X"99",X"d7",X"d7",X"d7",X"65",X"65",X"65",X"bd",
    X"99",X"99",X"d7",X"99",X"d7",X"99",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"bd",X"b4",X"01",X"01",
    X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",
    X"65",X"65",X"65",X"d7",X"65",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"bd",X"b4",X"b4",X"bd",X"bd",X"bd",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"65",X"65",X"65",X"d7",X"65",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",
    X"99",X"99",X"d7",X"99",X"d7",X"99",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"bd",X"b4",X"01",X"01",
    X"8a",X"8a",X"99",X"99",X"8a",X"99",X"99",X"99",X"99",X"d7",X"d7",X"d7",X"65",X"65",X"65",X"bd",
    X"2e",X"8a",X"8a",X"8a",X"2e",X"8a",X"8a",X"8a",X"99",X"99",X"99",X"d7",X"d7",X"65",X"bd",X"01",
    X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"99",X"99",X"d7",X"d7",X"65",X"bd",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"d7",X"65",X"bd",X"01",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",X"65",X"bd",X"bd",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"99",X"99",X"d7",X"65",X"bd",
    X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"8a",X"8a",X"99",X"99",X"d7",X"65",X"01",
    X"2e",X"8a",X"2e",X"2e",X"8a",X"8a",X"8a",X"8a",X"99",X"99",X"99",X"99",X"d7",X"d7",X"d7",X"65",
    X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"99",X"99",X"99",X"d7",X"d7",X"d7",X"65",X"65",X"bd",
    X"8a",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"bd",X"01",
    X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"65",X"bd",X"b4",X"01",X"01",
    X"65",X"65",X"d7",X"65",X"65",X"d7",X"65",X"65",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",
    X"b4",X"b4",X"65",X"bd",X"bd",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"65",X"65",X"d7",X"65",X"65",X"d7",X"65",X"65",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",
    X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"65",X"bd",X"b4",X"01",X"01",
    X"8a",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"bd",X"01",
    X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"99",X"99",X"99",X"d7",X"d7",X"d7",X"65",X"65",X"bd",
    X"2e",X"8a",X"2e",X"2e",X"8a",X"8a",X"8a",X"8a",X"99",X"99",X"99",X"99",X"d7",X"d7",X"d7",X"65",
    X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"8a",X"8a",X"99",X"99",X"d7",X"65",X"01",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"99",X"d7",X"d7",X"65",X"bd",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"99",X"d7",X"65",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",X"65",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"99",X"d7",X"bd",X"bd",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"65",X"bd",X"01",
    X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"99",X"99",X"d7",X"d7",X"65",X"bd",
    X"2e",X"8a",X"8a",X"8a",X"2e",X"8a",X"8a",X"8a",X"99",X"99",X"99",X"d7",X"d7",X"65",X"bd",X"01",
    X"8a",X"8a",X"99",X"99",X"8a",X"99",X"99",X"99",X"99",X"d7",X"d7",X"d7",X"65",X"65",X"65",X"bd",
    X"99",X"99",X"d7",X"99",X"d7",X"99",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"bd",X"b4",X"01",X"01",
    X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"65",X"65",X"65",X"bd",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"b4",X"bd",X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"99",X"99",X"d7",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"b4",X"65",X"d7",X"99",X"99",X"8a",X"99",X"99",X"d7",X"d7",X"65",X"01",X"01",
    X"01",X"01",X"65",X"bd",X"65",X"d7",X"99",X"8a",X"8a",X"8a",X"8a",X"99",X"d7",X"bd",X"01",X"01",
    X"01",X"01",X"d7",X"65",X"65",X"d7",X"d7",X"99",X"8a",X"99",X"99",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"65",X"d7",X"65",X"d7",X"99",X"8a",X"2e",X"8a",X"d7",X"d7",X"65",X"65",X"01",X"01",
    X"01",X"01",X"bd",X"65",X"d7",X"99",X"8a",X"8a",X"8a",X"8a",X"99",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"65",X"d7",X"d7",X"99",X"8a",X"99",X"99",X"d7",X"d7",X"65",X"65",X"01",X"01",
    X"01",X"01",X"01",X"65",X"65",X"d7",X"99",X"8a",X"8a",X"99",X"99",X"d7",X"65",X"d7",X"01",X"01",
    X"01",X"01",X"b4",X"65",X"d7",X"d7",X"d7",X"99",X"8a",X"8a",X"99",X"d7",X"d7",X"b4",X"01",X"01",
    X"01",X"01",X"bd",X"65",X"d7",X"d7",X"99",X"99",X"8a",X"99",X"99",X"d7",X"bd",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"b4",X"d7",X"99",X"99",X"8a",X"8a",X"99",X"d7",X"d7",X"bd",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"bd",X"65",X"d7",X"d7",X"99",X"99",X"d7",X"d7",X"65",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"65",X"bd",X"65",X"d7",X"99",X"8a",X"8a",X"99",X"99",X"d7",X"65",X"65",X"01",X"01",
    X"01",X"01",X"65",X"65",X"65",X"d7",X"99",X"8a",X"8a",X"99",X"d7",X"d7",X"65",X"d7",X"01",X"01",
    X"01",X"01",X"01",X"65",X"d7",X"99",X"99",X"8a",X"99",X"d7",X"d7",X"65",X"d7",X"65",X"01",X"01",
    X"01",X"01",X"01",X"65",X"d7",X"d7",X"99",X"8a",X"8a",X"99",X"d7",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"b4",X"bd",X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"8a",X"2e",X"8a",X"99",X"d7",X"bd",X"01",
    X"01",X"bd",X"b4",X"65",X"d7",X"99",X"99",X"8a",X"2e",X"8a",X"99",X"99",X"d7",X"d7",X"65",X"01",
    X"01",X"65",X"bd",X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"8a",X"8a",X"8a",X"99",X"d7",X"bd",X"01",
    X"01",X"d7",X"65",X"65",X"d7",X"d7",X"99",X"99",X"8a",X"99",X"99",X"99",X"d7",X"65",X"bd",X"01",
    X"01",X"65",X"d7",X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"8a",X"d7",X"d7",X"65",X"65",X"01",
    X"01",X"bd",X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",X"65",X"bd",X"01",
    X"01",X"bd",X"65",X"d7",X"d7",X"99",X"8a",X"8a",X"8a",X"99",X"99",X"d7",X"d7",X"65",X"65",X"01",
    X"01",X"01",X"65",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"65",X"d7",X"01",
    X"01",X"b4",X"65",X"d7",X"d7",X"d7",X"99",X"99",X"2e",X"8a",X"8a",X"99",X"d7",X"d7",X"b4",X"01",
    X"01",X"bd",X"65",X"d7",X"d7",X"99",X"99",X"8a",X"2e",X"8a",X"99",X"99",X"d7",X"bd",X"bd",X"01",
    X"01",X"bd",X"b4",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",X"bd",X"bd",X"01",
    X"01",X"bd",X"bd",X"65",X"d7",X"d7",X"99",X"8a",X"8a",X"99",X"d7",X"d7",X"65",X"65",X"bd",X"01",
    X"01",X"65",X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"65",X"65",X"01",
    X"01",X"65",X"65",X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"8a",X"99",X"d7",X"d7",X"65",X"d7",X"01",
    X"01",X"01",X"65",X"d7",X"99",X"99",X"8a",X"8a",X"8a",X"99",X"d7",X"d7",X"65",X"d7",X"65",X"01",
    X"01",X"01",X"65",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",X"65",X"bd",X"01",
    X"b4",X"01",X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"8a",X"2e",X"8a",X"99",X"d7",X"bd",
    X"bd",X"b4",X"65",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"d7",X"65",
    X"65",X"bd",X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"99",X"d7",X"bd",
    X"d7",X"65",X"65",X"d7",X"d7",X"d7",X"99",X"99",X"8a",X"8a",X"99",X"d7",X"99",X"d7",X"65",X"bd",
    X"65",X"d7",X"65",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"d7",X"d7",X"65",X"65",
    X"bd",X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",X"65",X"bd",
    X"bd",X"65",X"d7",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"d7",X"65",X"65",
    X"01",X"65",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"65",X"d7",
    X"b4",X"65",X"d7",X"d7",X"d7",X"d7",X"99",X"8a",X"8a",X"2e",X"8a",X"8a",X"99",X"d7",X"d7",X"b4",
    X"bd",X"65",X"d7",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"bd",X"bd",
    X"bd",X"b4",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",X"bd",X"bd",
    X"bd",X"bd",X"65",X"d7",X"d7",X"99",X"8a",X"2e",X"8a",X"8a",X"99",X"d7",X"d7",X"65",X"65",X"bd",
    X"65",X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"8a",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"65",X"65",
    X"65",X"65",X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"8a",X"2e",X"8a",X"99",X"d7",X"d7",X"65",X"d7",
    X"01",X"65",X"d7",X"99",X"99",X"8a",X"8a",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",X"65",X"d7",X"65",
    X"01",X"65",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",X"65",X"bd",
    X"65",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"65",X"bd",
    X"65",X"d7",X"99",X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",X"65",X"bd",
    X"bd",X"99",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"99",X"d7",X"65",
    X"b4",X"d7",X"99",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"8a",X"99",X"99",X"99",X"d7",X"65",X"65",
    X"bd",X"d7",X"d7",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"99",X"65",X"bd",
    X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"b4",
    X"bd",X"d7",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",X"65",X"b4",
    X"b4",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"65",X"bd",
    X"b4",X"d7",X"99",X"8a",X"8a",X"2e",X"8a",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",X"d7",X"65",X"bd",
    X"bd",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"d7",X"65",
    X"bd",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"65",
    X"65",X"65",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",X"65",X"b4",
    X"65",X"d7",X"99",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"8a",X"2e",X"8a",X"99",X"d7",X"65",X"bd",
    X"bd",X"d7",X"d7",X"99",X"8a",X"2e",X"8a",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",X"65",X"65",
    X"b4",X"65",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"99",X"d7",X"65",
    X"b4",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"65",X"65",
    X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",
    X"d7",X"99",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",X"65",
    X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"8a",X"99",X"d7",X"d7",
    X"65",X"d7",X"99",X"8a",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",
    X"65",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",X"d7",X"65",
    X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",
    X"d7",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",
    X"d7",X"d7",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"8a",X"8a",X"99",X"d7",
    X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",
    X"d7",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"d7",
    X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",
    X"d7",X"99",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"d7",X"d7",
    X"d7",X"d7",X"99",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",X"99",X"d7",
    X"d7",X"99",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"99",
    X"d7",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"99",X"d7",
    X"d7",X"d7",X"99",X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"65",X"65",X"bd",X"bd",X"bd",X"b4",X"01",X"bd",X"bd",X"65",X"d7",X"65",X"01",X"bd",
    X"65",X"65",X"65",X"bd",X"bd",X"b4",X"65",X"65",X"65",X"65",X"65",X"d7",X"65",X"65",X"65",X"65",
    X"d7",X"d7",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"65",X"d7",X"d7",X"d7",X"d7",X"d7",X"65",X"d7",
    X"d7",X"99",X"d7",X"d7",X"d7",X"99",X"d7",X"d7",X"d7",X"d7",X"99",X"d7",X"99",X"99",X"d7",X"99",
    X"99",X"99",X"99",X"99",X"d7",X"99",X"99",X"d7",X"99",X"99",X"8a",X"99",X"99",X"8a",X"99",X"8a",
    X"8a",X"8a",X"8a",X"8a",X"99",X"8a",X"99",X"d7",X"8a",X"8a",X"8a",X"8a",X"8a",X"8a",X"99",X"8a",
    X"8a",X"99",X"8a",X"8a",X"99",X"8a",X"8a",X"8a",X"8a",X"99",X"8a",X"2e",X"99",X"8a",X"8a",X"8a",
    X"99",X"d7",X"99",X"99",X"d7",X"99",X"99",X"8a",X"99",X"99",X"8a",X"8a",X"d7",X"8a",X"99",X"2e",
    X"d7",X"d7",X"d7",X"99",X"d7",X"d7",X"99",X"99",X"99",X"d7",X"99",X"d7",X"99",X"99",X"d7",X"99",
    X"d7",X"65",X"d7",X"d7",X"65",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",
    X"65",X"d7",X"65",X"65",X"65",X"bd",X"bd",X"d7",X"65",X"65",X"65",X"65",X"65",X"d7",X"65",X"65",
    X"bd",X"65",X"d7",X"65",X"bd",X"bd",X"bd",X"b4",X"d7",X"65",X"bd",X"65",X"bd",X"b4",X"bd",X"bd",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"bd",X"65",X"d7",X"65",X"bd",X"bd",X"bd",X"b4",X"d7",X"65",X"bd",X"65",X"bd",X"bd",X"65",X"bd",
    X"65",X"d7",X"65",X"65",X"65",X"bd",X"bd",X"d7",X"65",X"65",X"65",X"65",X"65",X"d7",X"d7",X"d7",
    X"d7",X"65",X"d7",X"d7",X"65",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"99",X"d7",X"99",
    X"d7",X"d7",X"d7",X"99",X"d7",X"d7",X"99",X"99",X"99",X"d7",X"99",X"d7",X"99",X"8a",X"99",X"8a",
    X"99",X"d7",X"99",X"99",X"d7",X"99",X"99",X"8a",X"99",X"99",X"8a",X"8a",X"d7",X"8a",X"99",X"2e",
    X"8a",X"99",X"8a",X"8a",X"99",X"8a",X"8a",X"8a",X"8a",X"99",X"8a",X"2e",X"99",X"8a",X"8a",X"8a",
    X"2e",X"8a",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",
    X"2e",X"8a",X"8a",X"2e",X"8a",X"2e",X"8a",X"99",X"2e",X"8a",X"2e",X"8a",X"99",X"8a",X"8a",X"8a",
    X"8a",X"8a",X"8a",X"8a",X"99",X"8a",X"99",X"d7",X"8a",X"8a",X"8a",X"99",X"d7",X"8a",X"99",X"99",
    X"99",X"99",X"99",X"99",X"d7",X"99",X"99",X"d7",X"99",X"99",X"8a",X"99",X"d7",X"99",X"99",X"d7",
    X"d7",X"99",X"d7",X"d7",X"d7",X"99",X"d7",X"d7",X"d7",X"d7",X"99",X"d7",X"d7",X"d7",X"d7",X"d7",
    X"d7",X"d7",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"65",X"d7",X"d7",X"65",X"65",X"65",X"65",X"65",
    X"65",X"65",X"65",X"bd",X"bd",X"b4",X"65",X"65",X"65",X"65",X"65",X"d7",X"65",X"bd",X"b4",X"01",
    X"01",X"01",X"65",X"65",X"bd",X"bd",X"bd",X"b4",X"01",X"bd",X"bd",X"65",X"d7",X"65",X"bd",X"b4",
    X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
    X"01",X"01",X"65",X"65",X"bd",X"bd",X"bd",X"b4",X"01",X"bd",X"bd",X"65",X"d7",X"65",X"bd",X"b4",
    X"65",X"65",X"65",X"bd",X"bd",X"b4",X"65",X"65",X"65",X"65",X"65",X"d7",X"65",X"bd",X"b4",X"01",
    X"d7",X"d7",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"65",X"d7",X"d7",X"65",X"65",X"65",X"65",X"65",
    X"d7",X"99",X"d7",X"d7",X"d7",X"99",X"d7",X"d7",X"d7",X"d7",X"99",X"d7",X"d7",X"d7",X"d7",X"d7",
    X"99",X"99",X"99",X"99",X"d7",X"99",X"99",X"d7",X"99",X"99",X"8a",X"99",X"d7",X"99",X"99",X"d7",
    X"8a",X"8a",X"8a",X"8a",X"99",X"8a",X"99",X"d7",X"8a",X"8a",X"8a",X"99",X"d7",X"8a",X"99",X"99",
    X"2e",X"8a",X"8a",X"2e",X"8a",X"2e",X"8a",X"99",X"2e",X"8a",X"2e",X"8a",X"99",X"8a",X"8a",X"8a",
    X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"99",X"2e",X"2e",X"8a",
    X"2e",X"2e",X"8a",X"2e",X"8a",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",
    X"2e",X"8a",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"8a",X"2e",X"8a",X"2e",
    X"8a",X"99",X"8a",X"8a",X"99",X"8a",X"8a",X"8a",X"8a",X"99",X"8a",X"2e",X"99",X"8a",X"8a",X"8a",
    X"99",X"d7",X"99",X"99",X"d7",X"99",X"99",X"8a",X"99",X"99",X"8a",X"8a",X"d7",X"8a",X"99",X"2e",
    X"d7",X"d7",X"d7",X"99",X"d7",X"d7",X"99",X"99",X"99",X"d7",X"99",X"d7",X"99",X"8a",X"99",X"8a",
    X"d7",X"65",X"d7",X"d7",X"65",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"99",X"d7",X"99",
    X"65",X"d7",X"65",X"65",X"65",X"bd",X"bd",X"d7",X"65",X"65",X"65",X"65",X"65",X"d7",X"d7",X"d7",
    X"bd",X"65",X"d7",X"65",X"bd",X"bd",X"bd",X"b4",X"d7",X"65",X"bd",X"65",X"bd",X"bd",X"65",X"bd",
    X"65",X"d7",X"65",X"65",X"65",X"bd",X"bd",X"d7",X"65",X"65",X"65",X"65",X"65",X"d7",X"d7",X"d7",
    X"d7",X"65",X"d7",X"d7",X"65",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"99",X"d7",X"99",
    X"d7",X"d7",X"d7",X"99",X"d7",X"d7",X"99",X"99",X"99",X"d7",X"99",X"d7",X"99",X"8a",X"99",X"8a",
    X"99",X"d7",X"99",X"99",X"d7",X"99",X"99",X"8a",X"99",X"99",X"8a",X"8a",X"d7",X"8a",X"99",X"2e",
    X"8a",X"99",X"8a",X"8a",X"99",X"8a",X"8a",X"8a",X"8a",X"99",X"8a",X"2e",X"99",X"8a",X"8a",X"8a",
    X"2e",X"8a",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"8a",X"2e",X"8a",X"2e",
    X"2e",X"2e",X"8a",X"2e",X"8a",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"99",X"2e",X"2e",X"8a",
    X"2e",X"8a",X"8a",X"2e",X"8a",X"2e",X"8a",X"99",X"2e",X"8a",X"2e",X"8a",X"99",X"8a",X"8a",X"8a",
    X"8a",X"8a",X"8a",X"8a",X"99",X"8a",X"99",X"d7",X"8a",X"8a",X"8a",X"99",X"d7",X"8a",X"99",X"99",
    X"99",X"99",X"99",X"99",X"d7",X"99",X"99",X"d7",X"99",X"99",X"8a",X"99",X"d7",X"99",X"99",X"d7",
    X"d7",X"99",X"d7",X"d7",X"d7",X"99",X"d7",X"d7",X"d7",X"d7",X"99",X"d7",X"d7",X"d7",X"d7",X"d7",
    X"d7",X"d7",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"65",X"d7",X"d7",X"65",X"65",X"65",X"65",X"65",
    X"65",X"65",X"65",X"bd",X"bd",X"b4",X"65",X"65",X"65",X"65",X"65",X"d7",X"65",X"bd",X"b4",X"01",
    X"d7",X"d7",X"65",X"65",X"65",X"d7",X"d7",X"d7",X"65",X"d7",X"d7",X"65",X"65",X"65",X"d7",X"d7",
    X"d7",X"99",X"d7",X"d7",X"d7",X"99",X"d7",X"d7",X"d7",X"d7",X"99",X"d7",X"d7",X"d7",X"d7",X"99",
    X"99",X"99",X"99",X"99",X"d7",X"99",X"99",X"d7",X"99",X"99",X"8a",X"99",X"d7",X"99",X"99",X"99",
    X"8a",X"8a",X"8a",X"8a",X"99",X"8a",X"99",X"d7",X"8a",X"8a",X"8a",X"99",X"d7",X"8a",X"99",X"8a",
    X"2e",X"8a",X"8a",X"2e",X"8a",X"2e",X"8a",X"99",X"2e",X"8a",X"2e",X"8a",X"99",X"8a",X"8a",X"8a",
    X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"99",X"2e",X"2e",X"8a",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"8a",X"2e",X"8a",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",
    X"2e",X"8a",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"8a",X"2e",X"8a",X"2e",
    X"8a",X"99",X"8a",X"8a",X"99",X"8a",X"8a",X"8a",X"8a",X"99",X"8a",X"2e",X"8a",X"8a",X"8a",X"8a",
    X"99",X"d7",X"99",X"99",X"d7",X"99",X"99",X"8a",X"99",X"99",X"8a",X"8a",X"99",X"8a",X"99",X"99",
    X"d7",X"d7",X"d7",X"99",X"d7",X"d7",X"99",X"99",X"99",X"d7",X"99",X"d7",X"99",X"99",X"d7",X"d7",
    X"d7",X"65",X"d7",X"d7",X"65",X"d7",X"d7",X"d7",X"d7",X"65",X"d7",X"65",X"d7",X"d7",X"d7",X"d7",
    X"01",X"01",X"b4",X"bd",X"65",X"65",X"d7",X"99",X"8a",X"8a",X"99",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"bd",X"65",X"65",X"d7",X"99",X"8a",X"2e",X"8a",X"99",X"d7",X"65",X"bd",X"01",X"01",
    X"bd",X"b4",X"bd",X"bd",X"65",X"d7",X"99",X"8a",X"8a",X"8a",X"8a",X"99",X"d7",X"65",X"b4",X"bd",
    X"bd",X"65",X"65",X"65",X"d7",X"d7",X"8a",X"8a",X"2e",X"8a",X"99",X"d7",X"d7",X"65",X"65",X"bd",
    X"d7",X"d7",X"d7",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",X"d7",X"d7",X"d7",
    X"99",X"d7",X"99",X"99",X"99",X"8a",X"8a",X"8a",X"2e",X"2e",X"8a",X"8a",X"99",X"99",X"d7",X"99",
    X"8a",X"99",X"8a",X"99",X"8a",X"99",X"8a",X"2e",X"2e",X"8a",X"2e",X"8a",X"99",X"8a",X"99",X"8a",
    X"2e",X"8a",X"8a",X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"2e",
    X"8a",X"8a",X"2e",X"2e",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"8a",X"8a",
    X"8a",X"8a",X"8a",X"99",X"8a",X"99",X"8a",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"8a",X"8a",X"8a",
    X"d7",X"99",X"99",X"d7",X"99",X"d7",X"99",X"8a",X"8a",X"2e",X"8a",X"99",X"d7",X"99",X"99",X"d7",
    X"d7",X"d7",X"d7",X"d7",X"d7",X"99",X"99",X"2e",X"8a",X"8a",X"99",X"d7",X"99",X"d7",X"d7",X"d7",
    X"bd",X"65",X"65",X"65",X"d7",X"d7",X"99",X"99",X"8a",X"8a",X"8a",X"d7",X"d7",X"65",X"65",X"bd",
    X"bd",X"b4",X"bd",X"65",X"65",X"d7",X"8a",X"8a",X"2e",X"8a",X"99",X"d7",X"65",X"bd",X"b4",X"bd",
    X"01",X"01",X"bd",X"bd",X"65",X"d7",X"99",X"2e",X"2e",X"8a",X"99",X"d7",X"65",X"bd",X"01",X"01",
    X"01",X"01",X"b4",X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"8a",X"d7",X"65",X"b4",X"01",X"01",
    X"01",X"01",X"bd",X"65",X"d7",X"d7",X"99",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",X"65",X"01",
    X"bd",X"bd",X"65",X"d7",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"65",X"bd",
    X"d7",X"65",X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"d7",
    X"99",X"d7",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"99",X"99",
    X"8a",X"99",X"99",X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"99",X"8a",X"99",
    X"8a",X"8a",X"8a",X"8a",X"8a",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"8a",
    X"8a",X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"8a",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",
    X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"8a",
    X"8a",X"8a",X"2e",X"8a",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"8a",X"8a",X"2e",X"8a",X"8a",X"8a",
    X"99",X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"8a",X"99",X"99",
    X"d7",X"99",X"99",X"8a",X"8a",X"2e",X"2e",X"8a",X"2e",X"8a",X"2e",X"2e",X"8a",X"2e",X"99",X"d7",
    X"d7",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"65",
    X"bd",X"65",X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"65",X"bd",
    X"bd",X"01",X"65",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"65",X"bd",X"bd",
    X"01",X"01",X"bd",X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"8a",X"99",X"d7",X"65",X"bd",X"01",
    X"01",X"bd",X"65",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"65",X"01",
    X"bd",X"65",X"d7",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",X"65",
    X"65",X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"d7",
    X"d7",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"8a",X"8a",X"99",X"d7",
    X"99",X"99",X"8a",X"8a",X"2e",X"99",X"99",X"8a",X"2e",X"2e",X"99",X"99",X"2e",X"8a",X"8a",X"99",
    X"8a",X"8a",X"2e",X"2e",X"8a",X"99",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"2e",X"8a",X"8a",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"8a",X"2e",X"8a",
    X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",
    X"8a",X"2e",X"2e",X"8a",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"2e",X"8a",X"8a",X"2e",X"2e",X"99",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"99",X"2e",X"2e",X"8a",
    X"99",X"8a",X"99",X"8a",X"2e",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"2e",X"2e",X"8a",
    X"99",X"99",X"8a",X"99",X"8a",X"2e",X"8a",X"2e",X"8a",X"2e",X"2e",X"2e",X"8a",X"8a",X"8a",X"8a",
    X"d7",X"d7",X"99",X"99",X"99",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"2e",X"8a",X"99",X"99",
    X"65",X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"8a",X"99",X"2e",X"8a",X"99",X"99",X"d7",
    X"bd",X"bd",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",X"65",
    X"01",X"bd",X"65",X"d7",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"65",X"01",
    X"65",X"d7",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"d7",X"65",X"bd",
    X"d7",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"99",X"d7",
    X"99",X"99",X"8a",X"8a",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"99",
    X"8a",X"8a",X"8a",X"2e",X"8a",X"99",X"99",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",
    X"2e",X"8a",X"2e",X"2e",X"2e",X"99",X"8a",X"8a",X"2e",X"2e",X"99",X"99",X"2e",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"99",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",
    X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"99",X"2e",X"2e",X"2e",X"8a",
    X"8a",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"2e",X"2e",X"8a",X"8a",
    X"99",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",
    X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",
    X"d7",X"d7",X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",X"65",
    X"65",X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"d7",X"65",X"bd",
    X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"8a",X"99",X"d7",
    X"99",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",
    X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",
    X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"99",X"2e",X"2e",X"8a",X"99",X"99",X"2e",X"2e",X"2e",X"8a",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"99",X"8a",X"99",X"2e",X"8a",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"8a",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"99",X"2e",X"2e",X"99",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"99",X"8a",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"8a",X"2e",X"2e",X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"2e",X"2e",X"2e",
    X"2e",X"2e",X"2e",X"2e",X"2e",X"99",X"99",X"2e",X"2e",X"2e",X"8a",X"99",X"99",X"2e",X"2e",X"2e",
    X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"99",X"2e",X"2e",X"8a",X"99",X"99",X"2e",X"2e",X"8a",X"8a",
    X"99",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",
    X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"99",X"99",
    X"d7",X"99",X"8a",X"8a",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"8a",X"8a",X"99",X"d7",others=>X"01"
    );
end package;