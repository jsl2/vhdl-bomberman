package touch_pkg is   
    type button_state is (none, up, right, down, left, bomb);
end;