use work.graphics_pkg.all;

package walls_pkg is    
    type walls_rom_type is array(0 to (2**11 - 1)) of pixel_type;    
    
    constant WALLS_FRAMES : walls_rom_type := 
   (X"00",X"fd",X"c4",X"29",X"c5",X"fd",X"c4",X"29",X"29",X"c4",X"c5",X"fd",X"c4",X"29",X"c5",X"fd",
    X"00",X"1f",X"af",X"af",X"29",X"1f",X"af",X"af",X"af",X"af",X"29",X"1f",X"af",X"af",X"29",X"1f",
    X"00",X"1f",X"82",X"82",X"c4",X"1f",X"82",X"82",X"82",X"82",X"29",X"1f",X"82",X"82",X"c4",X"1f",
    X"00",X"2e",X"82",X"2e",X"29",X"2e",X"82",X"b7",X"2e",X"b7",X"c4",X"2e",X"82",X"2e",X"29",X"2e",
    X"00",X"8f",X"82",X"82",X"c5",X"8f",X"82",X"82",X"82",X"82",X"c5",X"8f",X"82",X"82",X"b4",X"8f",
    X"00",X"1f",X"af",X"af",X"c5",X"1f",X"af",X"af",X"af",X"af",X"c5",X"1f",X"af",X"af",X"c5",X"1f",
    X"00",X"1f",X"af",X"af",X"c5",X"1f",X"af",X"af",X"af",X"af",X"c5",X"1f",X"af",X"af",X"c5",X"1f",
    X"00",X"1f",X"dc",X"83",X"c5",X"1f",X"83",X"c5",X"c5",X"c5",X"c5",X"1f",X"c5",X"c5",X"dc",X"1f",
    X"00",X"8f",X"8f",X"8f",X"8f",X"8f",X"8f",X"8f",X"8f",X"8f",X"8f",X"8f",X"8f",X"8f",X"8f",X"8f",
    X"00",X"fd",X"fd",X"fd",X"fd",X"fd",X"fd",X"3e",X"fd",X"fd",X"fd",X"fd",X"3e",X"fd",X"fd",X"3e",
    X"00",X"dc",X"dc",X"dc",X"dc",X"78",X"dc",X"dc",X"dc",X"dc",X"dc",X"dc",X"dc",X"dc",X"dc",X"1f",
    X"00",X"dc",X"00",X"00",X"dc",X"00",X"00",X"dc",X"8f",X"dc",X"3c",X"3c",X"dc",X"3c",X"00",X"1f",
    X"00",X"fd",X"83",X"00",X"fd",X"83",X"c5",X"00",X"3c",X"3c",X"83",X"00",X"fd",X"83",X"c5",X"1f",
    X"00",X"fd",X"96",X"c5",X"c5",X"c5",X"c5",X"c5",X"c5",X"c5",X"c5",X"c5",X"c5",X"96",X"c5",X"dc",
    X"00",X"fd",X"fd",X"fd",X"fd",X"fd",X"fd",X"fd",X"fd",X"fd",X"fd",X"fd",X"fd",X"fd",X"fd",X"fd",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"65",X"65",X"65",X"00",X"65",X"65",X"65",X"65",X"65",X"00",X"65",X"65",X"65",X"00",X"65",X"f9",
    X"bd",X"d7",X"d7",X"65",X"bd",X"d7",X"d7",X"d7",X"d7",X"65",X"bd",X"d7",X"d7",X"65",X"bd",X"f9",
    X"bd",X"99",X"99",X"65",X"bd",X"99",X"99",X"99",X"99",X"65",X"bd",X"99",X"99",X"65",X"bd",X"f9",
    X"2e",X"99",X"2e",X"65",X"2e",X"99",X"8a",X"2e",X"8a",X"65",X"2e",X"99",X"2e",X"65",X"2e",X"f9",
    X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"d7",X"99",X"f9",
    X"bd",X"d7",X"d7",X"00",X"bd",X"d7",X"d7",X"d7",X"d7",X"00",X"bd",X"d7",X"d7",X"d7",X"bd",X"f9",
    X"bd",X"d7",X"d7",X"00",X"bd",X"d7",X"d7",X"d7",X"d7",X"00",X"bd",X"d7",X"d7",X"d7",X"bd",X"f9",
    X"bd",X"65",X"00",X"00",X"bd",X"00",X"00",X"00",X"00",X"00",X"bd",X"00",X"00",X"65",X"bd",X"f9",
    X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"f9",
    X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"f9",
    X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"d7",X"f9",
    X"65",X"b4",X"65",X"00",X"65",X"65",X"d7",X"2e",X"65",X"00",X"65",X"b4",X"65",X"00",X"d7",X"f9",
    X"65",X"b4",X"65",X"00",X"65",X"b4",X"b4",X"b4",X"b4",X"00",X"65",X"b4",X"65",X"00",X"d7",X"f9",
    X"65",X"d7",X"b4",X"00",X"65",X"b4",X"d7",X"d7",X"65",X"00",X"65",X"b4",X"b4",X"d7",X"d7",X"f9",
    X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"f9",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"f9",
    X"65",X"65",X"65",X"00",X"65",X"65",X"65",X"65",X"65",X"00",X"65",X"65",X"65",X"00",X"65",X"f9",
    X"bd",X"99",X"99",X"65",X"bd",X"99",X"99",X"99",X"99",X"65",X"bd",X"99",X"99",X"65",X"bd",X"f9",
    X"2e",X"99",X"2e",X"65",X"2e",X"99",X"8a",X"2e",X"8a",X"65",X"2e",X"99",X"2e",X"65",X"2e",X"f9",
    X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"0f",X"99",X"f9",
    X"bd",X"d7",X"d7",X"0f",X"bd",X"0f",X"d7",X"d7",X"d7",X"00",X"bd",X"d7",X"d7",X"34",X"bd",X"f9",
    X"bd",X"d7",X"d7",X"00",X"bd",X"d7",X"d7",X"d7",X"d7",X"34",X"bd",X"d7",X"d7",X"d7",X"bd",X"f9",
    X"bd",X"65",X"00",X"00",X"bd",X"00",X"34",X"00",X"0f",X"00",X"bd",X"00",X"00",X"65",X"bd",X"f9",
    X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"34",X"99",X"99",X"99",X"34",X"99",X"99",X"f9",
    X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"34",X"f9",
    X"0f",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"0f",X"34",X"f9",
    X"65",X"65",X"0f",X"0f",X"34",X"65",X"34",X"65",X"65",X"65",X"0f",X"65",X"65",X"65",X"65",X"f9",
    X"65",X"b4",X"65",X"0f",X"65",X"65",X"d7",X"2e",X"65",X"00",X"65",X"0f",X"34",X"34",X"d7",X"f9",
    X"65",X"b4",X"65",X"00",X"65",X"b4",X"b4",X"34",X"b4",X"00",X"65",X"b4",X"65",X"0f",X"d7",X"f9",
    X"65",X"d7",X"b4",X"00",X"65",X"b4",X"d7",X"d7",X"65",X"00",X"65",X"b4",X"b4",X"d7",X"d7",X"f9",
    X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"f9",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"f9",
    X"65",X"65",X"65",X"00",X"65",X"65",X"65",X"65",X"65",X"00",X"65",X"65",X"65",X"00",X"65",X"f9",
    X"bd",X"99",X"0f",X"65",X"bd",X"99",X"99",X"99",X"99",X"65",X"bd",X"99",X"99",X"65",X"bd",X"f9",
    X"2e",X"99",X"34",X"65",X"2e",X"0f",X"8a",X"34",X"0f",X"65",X"2e",X"99",X"2e",X"65",X"2e",X"f9",
    X"99",X"99",X"34",X"00",X"99",X"34",X"99",X"34",X"34",X"00",X"99",X"99",X"34",X"0f",X"99",X"f9",
    X"bd",X"d7",X"d7",X"0f",X"bd",X"0f",X"34",X"d7",X"d7",X"00",X"bd",X"d7",X"34",X"34",X"bd",X"f9",
    X"bd",X"d7",X"0f",X"00",X"34",X"d7",X"d7",X"34",X"d7",X"34",X"bd",X"d7",X"0f",X"d7",X"bd",X"f9",
    X"bd",X"65",X"00",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"00",X"bd",X"00",X"00",X"0f",X"bd",X"f9",
    X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"34",X"f9",
    X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"34",X"f9",
    X"0f",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"0f",X"34",X"f9",
    X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"34",X"34",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"f9",
    X"65",X"b4",X"65",X"0f",X"0f",X"0f",X"d7",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"f9",
    X"65",X"b4",X"65",X"00",X"65",X"34",X"b4",X"34",X"b4",X"0f",X"65",X"b4",X"65",X"0f",X"d7",X"f9",
    X"65",X"d7",X"b4",X"00",X"65",X"b4",X"d7",X"d7",X"65",X"00",X"34",X"b4",X"b4",X"0f",X"d7",X"f9",
    X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"f9",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"f9",
    X"65",X"65",X"65",X"00",X"65",X"65",X"65",X"65",X"65",X"00",X"65",X"65",X"65",X"00",X"65",X"f9",
    X"bd",X"99",X"0f",X"65",X"bd",X"99",X"99",X"99",X"99",X"34",X"bd",X"99",X"99",X"65",X"bd",X"f9",
    X"2e",X"99",X"34",X"65",X"2e",X"0f",X"8a",X"34",X"0f",X"65",X"2e",X"34",X"2e",X"65",X"2e",X"f9",
    X"99",X"99",X"34",X"00",X"99",X"34",X"99",X"34",X"34",X"00",X"0f",X"99",X"34",X"0f",X"0f",X"f9",
    X"34",X"d7",X"0f",X"0f",X"bd",X"0f",X"34",X"34",X"0f",X"00",X"0f",X"d7",X"34",X"34",X"bd",X"f9",
    X"34",X"0f",X"0f",X"00",X"34",X"0f",X"d7",X"34",X"d7",X"34",X"bd",X"0f",X"0f",X"d7",X"bd",X"f9",
    X"0f",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"0f",X"34",X"f9",
    X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"34",X"f9",
    X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"34",X"f9",
    X"0f",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"0f",X"34",X"f9",
    X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"34",X"34",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"f9",
    X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"f9",
    X"65",X"b4",X"34",X"00",X"65",X"34",X"34",X"34",X"b4",X"0f",X"65",X"b4",X"65",X"0f",X"d7",X"f9",
    X"65",X"d7",X"34",X"00",X"0f",X"0f",X"34",X"d7",X"65",X"0f",X"34",X"b4",X"b4",X"0f",X"0f",X"f9",
    X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"f9",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"f9",
    X"65",X"65",X"65",X"00",X"65",X"65",X"65",X"65",X"65",X"00",X"65",X"0f",X"65",X"00",X"65",X"f9",
    X"bd",X"99",X"0f",X"65",X"bd",X"99",X"0f",X"99",X"99",X"34",X"bd",X"0f",X"0f",X"65",X"bd",X"f9",
    X"2e",X"0f",X"34",X"34",X"0f",X"0f",X"8a",X"34",X"0f",X"65",X"34",X"34",X"2e",X"0f",X"2e",X"f9",
    X"99",X"99",X"34",X"0f",X"99",X"34",X"34",X"34",X"34",X"0f",X"0f",X"99",X"34",X"0f",X"0f",X"f9",
    X"34",X"d7",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"00",X"0f",X"0f",X"34",X"34",X"0f",X"f9",
    X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"34",X"34",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"f9",
    X"0f",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"0f",X"34",X"f9",
    X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"34",X"f9",
    X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"34",X"f9",
    X"0f",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"0f",X"34",X"f9",
    X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"34",X"34",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"f9",
    X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"f9",
    X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"f9",
    X"0f",X"d7",X"34",X"00",X"0f",X"0f",X"34",X"34",X"65",X"0f",X"34",X"b4",X"b4",X"0f",X"0f",X"f9",
    X"b4",X"65",X"0f",X"65",X"b4",X"65",X"b4",X"65",X"b4",X"65",X"34",X"65",X"b4",X"65",X"b4",X"f9",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"f9",
    X"34",X"0f",X"65",X"0f",X"65",X"34",X"34",X"65",X"65",X"00",X"65",X"0f",X"65",X"00",X"65",X"f9",
    X"bd",X"99",X"0f",X"34",X"bd",X"99",X"0f",X"99",X"99",X"34",X"34",X"0f",X"0f",X"65",X"bd",X"f9",
    X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"65",X"34",X"34",X"0f",X"0f",X"2e",X"f9",
    X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"f9",
    X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"f9",
    X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"34",X"34",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"f9",
    X"0f",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"0f",X"34",X"f9",
    X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"34",X"f9",
    X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"34",X"0f",X"34",X"f9",
    X"0f",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"0f",X"34",X"f9",
    X"34",X"0f",X"0f",X"0f",X"34",X"0f",X"34",X"34",X"0f",X"34",X"0f",X"0f",X"0f",X"34",X"34",X"f9",
    X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"0f",X"34",X"34",X"0f",X"f9",
    X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"f9",
    X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"34",X"34",X"0f",X"0f",X"0f",X"f9",
    X"34",X"0f",X"0f",X"34",X"b4",X"65",X"b4",X"0f",X"b4",X"65",X"34",X"65",X"b4",X"34",X"b4",X"f9",
    X"34",X"0f",X"00",X"00",X"34",X"00",X"34",X"00",X"34",X"00",X"0f",X"0f",X"0f",X"00",X"0f",X"f9", others => X"01"
    );
end package;