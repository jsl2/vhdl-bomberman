library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package background_pkg is
    type bg_rom_type is array(0 to (2**17 - 1)) of std_logic_vector(7 downto 0);
    constant BG_PIC : bg_rom_type := (X"0b",X"33",X"f0",X"6d",X"3f",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"54",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"54",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"54",X"1a",X"6d",X"3f",X"98",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"0d",X"54",X"1a",X"6d",X"3f",X"54",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"54",X"1a",X"6d",X"3f",X"54",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"54",X"1a",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"17",X"0b",X"61",X"33",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"54",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"54",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"54",X"1a",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"98",X"0b",
    X"98",X"17",X"84",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"3f",X"6d",X"f0",X"6d",X"3f",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"61",X"ad",X"6d",X"f0",X"17",X"98",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"3f",X"54",X"98",X"3b",X"17",
    X"aa",X"ba",X"17",X"98",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"6d",X"f0",X"6d",X"f0",X"6d",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"2c",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"2c",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"79",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"98",X"1b",X"33",X"f0",X"12",X"98",X"3b",X"98",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"3f",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"6d",X"61",X"ad",X"98",X"3f",
    X"aa",X"7c",X"61",X"3b",X"98",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"1a",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"2c",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"79",X"6d",X"f0",X"6d",X"79",X"6d",X"f0",X"6d",X"f0",X"6d",X"79",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"79",X"6d",X"f0",X"6d",X"f0",X"6d",X"79",X"6d",X"6d",X"f0",X"6d",X"79",X"6d",X"f0",X"6d",X"6d",X"f0",X"6d",X"1a",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"79",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"79",X"6d",X"f0",X"6d",X"79",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"79",X"6d",X"f0",X"6d",X"79",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"79",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"98",X"3b",X"98",X"6d",X"6d",X"aa",X"aa",X"6d",X"3b",X"98",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"1a",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"33",X"17",X"98",X"f0",X"6d",
    X"9e",X"aa",X"7c",X"61",X"58",X"33",X"3b",X"33",X"33",X"3b",X"33",X"33",X"53",X"33",X"33",X"3b",X"33",X"3b",X"33",X"33",X"33",X"3b",X"33",X"33",X"33",X"3b",X"33",X"33",X"33",X"33",X"3b",X"33",X"3b",X"33",X"53",X"33",X"33",X"33",X"3b",X"33",X"33",X"33",X"33",X"3b",X"33",X"3b",X"33",X"33",X"53",X"33",X"33",X"98",X"3b",X"33",X"98",X"33",X"53",X"33",X"33",X"53",X"33",X"33",X"33",X"33",X"3b",X"98",X"33",X"33",X"33",X"53",X"33",X"33",X"33",X"3b",X"33",X"33",X"33",X"53",X"33",X"3b",X"33",X"33",X"33",X"3b",X"33",X"33",X"3b",X"33",X"33",X"33",X"3b",X"61",X"33",X"33",X"3b",X"98",X"3b",X"33",X"33",X"33",X"3b",X"33",X"33",X"33",X"33",X"3b",X"33",X"33",X"3b",X"33",X"33",X"3b",X"33",X"33",X"3b",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"3b",X"33",X"33",X"33",X"33",X"3b",X"33",X"33",X"33",X"33",X"33",X"17",X"33",X"33",X"33",X"3b",X"33",X"3b",X"33",X"33",X"17",X"33",X"33",X"33",X"3b",X"33",X"3b",X"33",X"33",X"17",X"33",X"33",X"33",X"3b",X"33",X"3b",X"33",X"33",X"17",X"33",X"33",X"33",X"3b",X"33",X"3b",X"33",X"33",X"3b",X"33",X"33",X"33",X"cd",X"33",X"3b",X"33",X"33",X"17",X"33",X"33",X"33",X"3b",X"33",X"cd",X"33",X"33",X"17",X"33",X"33",X"33",X"3b",X"33",X"cd",X"33",X"33",X"3b",X"33",X"33",X"33",X"3b",X"33",X"3b",X"33",X"33",X"17",X"33",X"33",X"33",X"cd",X"33",X"3b",X"33",X"33",X"53",X"3b",X"33",X"33",X"17",X"53",X"33",X"3b",X"33",X"3b",X"33",X"3b",X"33",X"33",X"17",X"33",X"33",X"53",X"33",X"17",X"33",X"33",X"3b",X"33",X"3b",X"33",X"17",X"33",X"33",X"53",X"33",X"17",X"33",X"33",X"3b",X"33",X"cd",X"33",X"17",X"33",X"33",X"53",X"33",X"17",X"33",X"33",X"cd",X"33",X"3b",X"33",X"17",X"33",X"33",X"53",X"33",X"17",X"33",X"33",X"cd",X"33",X"3b",X"33",X"3b",X"33",X"33",X"53",X"33",X"17",X"33",X"33",X"cd",X"33",X"3b",X"33",X"17",X"33",X"33",X"53",X"33",X"17",X"33",X"33",X"3b",X"33",X"3b",X"33",X"17",X"33",X"33",X"53",X"33",X"17",X"33",X"33",X"3b",X"33",X"3b",X"33",X"17",X"33",X"33",X"53",X"33",X"17",X"33",X"33",X"3b",X"33",X"3b",X"33",X"17",X"33",X"33",X"53",X"33",X"17",X"33",X"33",X"cd",X"33",X"3b",X"33",X"17",X"33",X"33",X"53",X"33",X"17",X"33",X"33",X"3b",X"33",X"3b",X"33",X"17",X"33",X"cd",X"33",X"17",X"3b",X"98",X"f0",X"6d",X"f0",X"aa",X"60",X"aa",X"98",X"3b",X"84",X"33",X"3b",X"33",X"33",X"33",X"33",X"33",X"3b",X"33",X"33",X"33",X"33",X"53",X"33",X"33",X"3b",X"33",X"33",X"3b",X"33",X"33",X"33",X"3b",X"33",X"33",X"33",X"33",X"3b",X"33",X"33",X"33",X"33",X"3b",X"33",X"33",X"3b",X"33",X"33",X"33",X"3b",X"33",X"33",X"17",X"33",X"33",X"17",X"33",X"33",X"3b",X"33",X"53",X"33",X"3b",X"33",X"33",X"3b",X"33",X"3b",X"33",X"33",X"53",X"33",X"33",X"53",X"33",X"3b",X"33",X"53",X"33",X"3b",X"33",X"33",X"3b",X"33",X"3b",X"33",X"33",X"33",X"3b",X"33",X"33",X"53",X"33",X"3b",X"33",X"33",X"3b",X"33",X"33",X"3b",X"33",X"33",X"3b",X"33",X"33",X"3b",X"33",X"33",X"33",X"17",X"33",X"3b",X"33",X"3b",X"33",X"33",X"33",X"3b",X"98",X"17",X"98",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"0b",X"1b",X"83",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"83",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"83",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"83",X"e4",X"0b",X"0b",X"0b",X"83",X"0b",X"1b",X"0b",X"c5",X"1b",X"0b",X"0b",X"1b",X"c5",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"1b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"1b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"1b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"1b",X"83",X"0b",X"1b",X"0b",X"56",X"1b",X"0b",X"0b",X"1b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"1b",X"83",X"0b",X"1b",X"0b",X"56",X"1b",X"0b",X"0b",X"1b",X"56",X"0b",X"1b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"56",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"56",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"1b",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"3f",X"6d",X"42",X"6d",X"12",X"98",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"83",X"0b",X"3c",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"33",X"6d",X"3f",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"aa",X"84",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"ad",X"0b",X"1b",X"0b",X"0b",X"ad",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"ad",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"ad",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"e4",X"0b",X"0b",X"1b",X"0b",X"0b",X"e4",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"83",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"3c",X"0b",X"1b",X"0b",X"1b",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"3c",X"0b",X"1b",X"0b",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"0b",X"0b",X"3c",X"0b",X"1b",X"0b",X"3c",X"0b",X"1b",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"00",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"3b",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"60",X"aa",X"7c",X"61",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"ad",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"ad",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"ad",X"0b",X"0b",X"ad",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"ad",X"0b",X"0b",X"0b",X"ad",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"ad",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"ad",X"0b",X"1b",X"0b",X"1b",X"0b",X"e4",X"0b",X"e4",X"0b",X"e4",X"0b",X"e4",X"0b",X"e4",X"0b",X"e4",X"0b",X"e4",X"0b",X"e4",X"0b",X"e4",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"3c",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"5d",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"5d",X"0b",X"1b",X"0b",X"5d",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"5d",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"5d",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"3c",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"3c",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"3c",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"6d",X"aa",X"7c",X"9e",X"98",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"3c",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"83",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"3c",X"0b",X"1b",X"0b",X"3c",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"aa",X"9e",X"aa",X"84",X"0b",X"1b",X"0b",X"61",X"2f",X"2f",X"2f",X"f0",X"2f",X"2f",X"28",X"2f",X"2f",X"f0",X"79",X"2f",X"2f",X"2f",X"28",X"2f",X"2f",X"f0",X"2f",X"2f",X"2f",X"f0",X"2f",X"28",X"2f",X"28",X"2f",X"2f",X"f0",X"2f",X"f0",X"2f",X"2f",X"2f",X"69",X"2f",X"f0",X"2f",X"28",X"2f",X"2f",X"2f",X"2f",X"2f",X"28",X"2f",X"28",X"2f",X"79",X"2f",X"2f",X"28",X"2f",X"2f",X"f0",X"2f",X"2f",X"2f",X"28",X"2f",X"28",X"2f",X"f0",X"28",X"ed",X"79",X"2f",X"f0",X"2f",X"79",X"2f",X"28",X"2f",X"28",X"2f",X"2f",X"f0",X"2f",X"2f",X"2f",X"28",X"f0",X"f0",X"28",X"3f",X"12",X"63",X"69",X"69",X"16",X"4c",X"16",X"69",X"4c",X"16",X"12",X"3f",X"1a",X"f0",X"f0",X"2f",X"79",X"2f",X"2f",X"2f",X"28",X"2f",X"2f",X"f0",X"2f",X"2f",X"2f",X"f0",X"79",X"2f",X"2f",X"f0",X"ed",X"2f",X"f0",X"00",X"00",X"00",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"12",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"19",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"75",X"03",X"03",X"75",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"27",X"19",X"03",X"03",X"b2",X"19",X"03",X"03",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"03",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"b2",X"27",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"0b",X"3c",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"7c",X"aa",X"7c",X"61",X"0b",X"0b",X"0b",X"2f",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"75",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"2e",X"ec",X"03",X"1a",X"03",X"1a",X"03",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"b2",X"03",X"b2",X"03",X"75",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"03",X"14",X"09",X"ec",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"09",X"14",X"03",X"03",X"71",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"00",X"00",X"00",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"3b",X"6d",X"f0",X"3f",X"6d",X"aa",X"9e",X"aa",X"92",X"61",X"0b",X"0b",X"0b",X"03",X"1a",X"03",X"03",X"19",X"03",X"1a",X"03",X"03",X"19",X"b2",X"19",X"71",X"03",X"1a",X"71",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"71",X"19",X"b2",X"19",X"b2",X"27",X"19",X"03",X"b2",X"03",X"75",X"03",X"03",X"1a",X"03",X"19",X"b2",X"19",X"b2",X"03",X"b2",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"27",X"1a",X"03",X"19",X"03",X"0b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"1b",X"83",X"2f",X"19",X"b2",X"27",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"27",X"75",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"27",X"19",X"03",X"19",X"b2",X"03",X"2e",X"0b",X"2e",X"03",X"1a",X"03",X"03",X"19",X"b2",X"27",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"71",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"03",X"b2",X"03",X"03",X"03",X"14",X"68",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"14",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"b2",X"27",X"19",X"71",X"19",X"71",X"19",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"00",X"00",X"00",X"82",X"3c",X"82",X"3c",X"82",X"00",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"00",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"19",X"03",X"1a",X"03",X"b2",X"27",X"03",X"03",X"1a",X"b2",X"03",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"27",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"27",X"1b",X"0b",X"1b",X"17",X"f0",X"6d",X"3f",X"6d",
    X"aa",X"7c",X"0d",X"9e",X"98",X"0b",X"0b",X"1b",X"2f",X"03",X"03",X"b2",X"19",X"71",X"19",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"2e",X"00",X"1b",X"2e",X"03",X"b2",X"19",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"19",X"b2",X"27",X"19",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"14",X"14",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"14",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"f0",X"6d",X"6d",X"f0",X"60",X"aa",X"60",X"aa",X"98",X"0b",X"1b",X"0b",X"d8",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"03",X"75",X"03",X"03",X"b2",X"27",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"19",X"03",X"19",X"03",X"75",X"03",X"75",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"ad",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"7c",X"aa",X"61",X"0b",X"1b",X"0b",X"2f",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"71",X"19",X"03",X"1a",X"03",X"75",X"03",X"b2",X"d8",X"19",X"03",X"1a",X"03",X"19",X"03",X"03",X"03",X"2e",X"0b",X"0b",X"2e",X"03",X"19",X"03",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"19",X"71",X"03",X"14",X"14",X"09",X"68",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"14",X"03",X"03",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"19",X"03",X"b2",X"00",X"00",X"00",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"53",X"6d",X"f0",X"3f",X"6d",X"aa",X"aa",X"aa",X"9e",X"98",X"0b",X"0b",X"0b",X"03",X"1a",X"03",X"71",X"75",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"03",X"75",X"03",X"b2",X"03",X"03",X"19",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"75",X"03",X"0b",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"9e",X"aa",X"60",X"98",X"0b",X"0b",X"1b",X"2f",X"19",X"03",X"b2",X"03",X"b2",X"27",X"75",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"19",X"71",X"19",X"71",X"27",X"03",X"19",X"b2",X"03",X"b2",X"03",X"19",X"71",X"03",X"03",X"14",X"2e",X"1b",X"3c",X"2e",X"03",X"b2",X"03",X"b2",X"19",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"d8",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"03",X"14",X"14",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"68",X"14",X"03",X"03",X"19",X"b2",X"27",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"19",X"00",X"00",X"fb",X"f4",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"fb",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"7c",X"9e",X"aa",X"98",X"0b",X"1b",X"0b",X"19",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"19",X"b2",X"27",X"19",X"03",X"75",X"03",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"75",X"03",X"75",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"75",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"0b",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"79",X"03",X"b2",X"19",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"19",X"b2",X"27",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"03",X"03",X"14",X"2e",X"75",X"0b",X"2e",X"4d",X"19",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"19",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"03",X"03",X"14",X"09",X"ec",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"09",X"14",X"03",X"03",X"71",X"27",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"19",X"03",X"b2",X"00",X"00",X"f4",X"3c",X"00",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"4f",X"f4",X"00",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"9e",X"aa",X"aa",X"7c",X"61",X"0b",X"0b",X"1b",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"75",X"03",X"03",X"b2",X"19",X"03",X"75",X"03",X"1a",X"03",X"71",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"27",X"03",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"0b",X"3c",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"60",X"aa",X"92",X"61",X"0b",X"0b",X"83",X"2f",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"d8",X"14",X"09",X"2e",X"19",X"00",X"2e",X"4d",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"21",X"03",X"1a",X"03",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"71",X"27",X"19",X"03",X"b2",X"03",X"b2",X"03",X"03",X"14",X"68",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"14",X"27",X"d8",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"f4",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"fb",X"f4",X"fb",X"f4",X"f4",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",X"aa",X"7c",X"aa",X"9e",X"98",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"1a",X"03",X"03",X"b2",X"19",X"03",X"03",X"03",X"1a",X"03",X"19",X"71",X"19",X"71",X"19",X"71",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"71",X"19",X"71",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"1b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"2f",X"03",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"71",X"d8",X"14",X"09",X"2e",X"75",X"1b",X"25",X"ec",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"2e",X"2e",X"03",X"1a",X"03",X"b2",X"27",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"03",X"14",X"09",X"14",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"14",X"03",X"03",X"71",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"60",X"aa",X"12",X"aa",X"98",X"0b",X"0b",X"0b",X"19",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"75",X"03",X"03",X"1a",X"03",X"19",X"71",X"19",X"71",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"19",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"d8",X"19",X"03",X"b2",X"03",X"b2",X"27",X"19",X"03",X"19",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"03",X"71",X"19",X"03",X"19",X"03",X"b2",X"27",X"75",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"0b",X"0b",X"0b",X"3b",X"3f",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"60",X"61",X"0b",X"1b",X"0b",X"2f",X"19",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"03",X"03",X"14",X"68",X"14",X"2e",X"19",X"3c",X"25",X"ec",X"03",X"1a",X"ec",X"03",X"1a",X"03",X"03",X"cc",X"0b",X"2e",X"03",X"1a",X"03",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"14",X"09",X"68",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"14",X"14",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"d8",X"19",X"03",X"b2",X"d8",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"91",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"aa",X"2c",X"aa",X"84",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"75",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"71",X"19",X"71",X"03",X"1a",X"03",X"71",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"19",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"19",X"71",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"1b",X"0b",X"1b",X"98",X"6d",X"f0",X"3f",X"6d",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"0b",X"0b",X"79",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"75",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"03",X"03",X"14",X"09",X"09",X"2e",X"4d",X"1b",X"4d",X"2e",X"03",X"19",X"2e",X"2e",X"03",X"1a",X"03",X"2e",X"1b",X"75",X"2e",X"03",X"19",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"b2",X"d8",X"03",X"1a",X"03",X"1a",X"03",X"03",X"71",X"d8",X"03",X"14",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"14",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"d8",X"1a",X"03",X"b2",X"d8",X"19",X"71",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"3b",X"6d",X"f0",X"6d",X"f0",X"aa",X"12",X"aa",X"aa",X"98",X"0b",X"0b",X"0b",X"d8",X"1a",X"03",X"71",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"75",X"03",X"b2",X"03",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"75",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"27",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"19",X"03",X"19",X"0b",X"0b",X"0b",X"3b",X"f0",X"6d",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"60",X"98",X"1b",X"0b",X"1b",X"2f",X"03",X"75",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"1a",X"03",X"71",X"03",X"03",X"14",X"09",X"09",X"ec",X"2e",X"4d",X"1b",X"4d",X"2e",X"03",X"b2",X"2e",X"3c",X"2e",X"03",X"1a",X"ec",X"0b",X"75",X"2e",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"75",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"19",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"03",X"14",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"a7",X"03",X"03",X"03",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"19",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"4a",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"3f",X"6d",X"aa",X"7c",X"9e",X"98",X"1b",X"0b",X"1b",X"03",X"1a",X"03",X"75",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"71",X"19",X"71",X"27",X"19",X"03",X"1a",X"03",X"b2",X"27",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"71",X"19",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"1b",X"0b",X"1b",X"33",X"6d",X"f0",X"f0",X"6d",
    X"9e",X"aa",X"9e",X"aa",X"98",X"0b",X"0b",X"0b",X"79",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"d8",X"14",X"09",X"68",X"14",X"ec",X"e9",X"3c",X"75",X"2e",X"1a",X"03",X"cc",X"0b",X"75",X"2e",X"03",X"cc",X"0b",X"19",X"2e",X"03",X"2e",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"75",X"03",X"1a",X"03",X"71",X"19",X"71",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"27",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"14",X"ec",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"09",X"14",X"03",X"03",X"71",X"19",X"71",X"03",X"19",X"03",X"1a",X"03",X"b2",X"27",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"71",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"12",X"aa",X"aa",X"84",X"0b",X"0b",X"0b",X"19",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"b2",X"27",X"75",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"75",X"03",X"19",X"71",X"19",X"03",X"19",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"19",X"1a",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"71",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"6d",X"3f",
    X"aa",X"9e",X"7c",X"aa",X"84",X"0b",X"1b",X"0b",X"2f",X"19",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"71",X"d8",X"2e",X"09",X"09",X"ec",X"2e",X"25",X"3c",X"19",X"2e",X"03",X"03",X"2e",X"1b",X"19",X"2e",X"03",X"cc",X"1b",X"75",X"2e",X"19",X"ec",X"2e",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"71",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"19",X"71",X"19",X"03",X"03",X"b2",X"03",X"2e",X"03",X"03",X"03",X"14",X"09",X"68",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"09",X"14",X"03",X"03",X"03",X"75",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"d8",X"75",X"03",X"03",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"f4",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",X"42",X"6d",X"aa",X"7c",X"61",X"0b",X"1b",X"0b",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"19",X"71",X"19",X"71",X"19",X"03",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"75",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"19",X"71",X"19",X"03",X"71",X"27",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"1b",X"0b",X"1b",X"3b",X"6d",X"f0",X"3f",X"54",
    X"aa",X"7c",X"aa",X"aa",X"ba",X"0b",X"0b",X"0b",X"f0",X"03",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"27",X"75",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"03",X"2e",X"2e",X"09",X"09",X"4d",X"2e",X"1b",X"75",X"2e",X"03",X"1a",X"ec",X"0b",X"75",X"2e",X"03",X"cc",X"0b",X"19",X"2e",X"03",X"2e",X"0b",X"2e",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"d8",X"19",X"71",X"19",X"03",X"19",X"71",X"19",X"03",X"b2",X"27",X"03",X"21",X"03",X"1a",X"03",X"03",X"cc",X"2e",X"03",X"03",X"03",X"14",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"14",X"14",X"03",X"03",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"03",X"b2",X"03",X"03",X"19",X"b2",X"27",X"03",X"1a",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"70",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"6d",X"aa",X"9e",X"aa",X"98",X"0b",X"0b",X"0b",X"d8",X"1a",X"03",X"b2",X"27",X"19",X"71",X"19",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"19",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"19",X"b2",X"27",X"19",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"0b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"9e",X"aa",X"aa",X"60",X"98",X"0b",X"1b",X"0b",X"2f",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"71",X"03",X"2e",X"1b",X"2e",X"09",X"4d",X"2e",X"3c",X"75",X"2e",X"4d",X"03",X"2e",X"3c",X"75",X"2e",X"03",X"e5",X"3c",X"75",X"2e",X"ec",X"2e",X"1b",X"0b",X"2e",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"b2",X"27",X"19",X"71",X"19",X"71",X"19",X"03",X"b2",X"19",X"b2",X"19",X"2e",X"2e",X"03",X"1a",X"03",X"2e",X"1b",X"2e",X"03",X"03",X"14",X"14",X"09",X"2e",X"2e",X"2e",X"2e",X"09",X"14",X"03",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"19",X"03",X"75",X"03",X"b2",X"03",X"03",X"1a",X"03",X"00",X"00",X"fb",X"00",X"a4",X"91",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"79",X"6d",X"f0",X"6d",X"aa",X"aa",X"7c",X"9e",X"98",X"0b",X"1b",X"0b",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"19",X"71",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"03",X"1a",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"75",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"3c",X"0b",X"0b",X"3b",X"1a",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"9e",X"aa",X"98",X"0b",X"83",X"1b",X"ed",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"03",X"03",X"1a",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"71",X"19",X"03",X"03",X"1a",X"03",X"03",X"cc",X"0b",X"3c",X"2e",X"14",X"2e",X"1b",X"3c",X"2e",X"4d",X"19",X"21",X"0b",X"19",X"2e",X"03",X"cc",X"0b",X"75",X"2e",X"2e",X"2e",X"3c",X"1b",X"2e",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"03",X"03",X"2e",X"1b",X"2e",X"03",X"1a",X"2e",X"3c",X"0b",X"2e",X"03",X"14",X"09",X"09",X"ec",X"2e",X"2e",X"09",X"68",X"14",X"d8",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f4",X"4f",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"12",X"aa",X"aa",X"aa",X"98",X"0b",X"0b",X"3c",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"27",X"75",X"b2",X"03",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"75",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"71",X"19",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"75",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"d8",X"0b",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"77",X"03",X"1a",X"03",X"75",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"0b",X"1b",X"3c",X"0b",X"1b",X"3c",X"0b",X"3c",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"2e",X"00",X"0b",X"2e",X"2e",X"2e",X"0b",X"3c",X"25",X"ec",X"03",X"2e",X"1b",X"75",X"2e",X"03",X"cc",X"1b",X"3c",X"e9",X"30",X"2e",X"0b",X"1b",X"3d",X"2e",X"03",X"03",X"b2",X"d8",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"03",X"19",X"03",X"71",X"19",X"71",X"03",X"19",X"71",X"19",X"b2",X"2e",X"3c",X"0b",X"2e",X"03",X"30",X"1b",X"0b",X"2e",X"03",X"2e",X"14",X"09",X"2e",X"2e",X"2e",X"ec",X"14",X"14",X"03",X"71",X"27",X"19",X"03",X"1a",X"03",X"b2",X"03",X"75",X"03",X"1a",X"03",X"03",X"b2",X"27",X"75",X"03",X"03",X"b2",X"03",X"03",X"1a",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f4",X"2e",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"fb",X"f4",X"fb",X"f4",X"91",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"3b",X"6d",X"3f",X"6d",X"f0",X"aa",X"60",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"b2",X"03",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"71",X"27",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"d8",X"75",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"75",X"03",X"03",X"1a",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"b2",X"27",X"75",X"03",X"19",X"71",X"19",X"03",X"19",X"b2",X"cd",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"79",X"03",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"3c",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"0b",X"03",X"19",X"03",X"1a",X"03",X"03",X"71",X"2e",X"0b",X"3c",X"2e",X"2e",X"ec",X"75",X"1b",X"4d",X"2e",X"19",X"ec",X"0b",X"75",X"2e",X"03",X"e5",X"3c",X"0b",X"3d",X"2e",X"ec",X"75",X"0b",X"25",X"ec",X"03",X"1a",X"03",X"b2",X"27",X"75",X"03",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"2e",X"0b",X"00",X"2e",X"03",X"2e",X"0b",X"00",X"2e",X"03",X"2e",X"2e",X"14",X"2e",X"2e",X"2e",X"09",X"14",X"27",X"03",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"71",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"2e",X"fb",X"f4",X"fb",X"f4",X"91",X"f4",X"f4",X"fb",X"f4",X"3c",X"00",X"f4",X"fb",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"60",X"aa",X"36",X"aa",X"33",X"0b",X"0b",X"1b",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"19",X"b2",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"71",X"19",X"71",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"75",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"0b",X"0b",X"0b",X"17",X"6d",X"3f",X"6d",X"f0",
    X"9e",X"aa",X"9e",X"aa",X"98",X"0b",X"0b",X"0b",X"79",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"03",X"0b",X"00",X"2e",X"0b",X"3c",X"0b",X"0b",X"3c",X"03",X"b2",X"03",X"03",X"71",X"19",X"03",X"2e",X"1b",X"3c",X"e9",X"30",X"2e",X"19",X"0b",X"4d",X"2e",X"03",X"2e",X"0b",X"3c",X"2e",X"03",X"2e",X"0b",X"0b",X"4d",X"2e",X"2e",X"19",X"3c",X"4d",X"2e",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"75",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"19",X"71",X"27",X"03",X"1a",X"ec",X"0b",X"0b",X"2e",X"1a",X"2e",X"1b",X"0b",X"2e",X"ec",X"2e",X"0b",X"ec",X"09",X"2e",X"2e",X"2e",X"09",X"14",X"03",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"2e",X"2e",X"fb",X"f4",X"fb",X"f4",X"fb",X"91",X"f4",X"fb",X"f4",X"fb",X"00",X"fb",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"60",X"aa",X"98",X"1b",X"0b",X"0b",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"19",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"b2",X"27",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"75",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"0b",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"84",X"0b",X"0b",X"1b",X"ed",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"b2",X"03",X"0b",X"1b",X"2e",X"2e",X"3c",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"ec",X"bf",X"0b",X"3d",X"2e",X"2e",X"75",X"3c",X"75",X"2e",X"2e",X"2e",X"3c",X"0b",X"ec",X"2e",X"2e",X"3c",X"0b",X"4d",X"2e",X"ec",X"bf",X"0b",X"4d",X"2e",X"03",X"b2",X"03",X"19",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"75",X"03",X"1a",X"03",X"2e",X"00",X"1b",X"2e",X"03",X"cc",X"3c",X"0b",X"2e",X"2e",X"2e",X"1b",X"0b",X"2e",X"2e",X"2e",X"09",X"14",X"03",X"03",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"03",X"19",X"03",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"fb",X"00",X"2e",X"fb",X"f4",X"4f",X"f4",X"fb",X"f4",X"4f",X"f4",X"fb",X"f4",X"00",X"fb",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"53",X"6d",X"f0",X"3f",X"6d",X"aa",X"60",X"42",X"6d",X"ba",X"0b",X"0b",X"1b",X"03",X"b2",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"75",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"75",X"03",X"19",X"03",X"b2",X"03",X"75",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"03",X"1a",X"03",X"b2",X"27",X"75",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"0b",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"9e",X"aa",X"7c",X"61",X"0b",X"0b",X"0b",X"79",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"03",X"0b",X"0b",X"ec",X"1b",X"3c",X"0b",X"1b",X"0b",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"2e",X"75",X"1b",X"4d",X"2e",X"ec",X"19",X"0b",X"75",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"00",X"1b",X"19",X"2e",X"2e",X"4d",X"1b",X"75",X"2e",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"2e",X"0b",X"0b",X"2e",X"03",X"2e",X"0b",X"1b",X"2e",X"2e",X"2e",X"3c",X"0b",X"2e",X"2e",X"09",X"09",X"2e",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"19",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"2e",X"fb",X"00",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"2e",X"2e",X"fb",X"00",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"aa",X"6d",X"aa",X"74",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"27",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"19",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"1b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"0d",X"9e",X"98",X"0b",X"1b",X"0b",X"2f",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"03",X"b2",X"1b",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"0b",X"27",X"19",X"03",X"b2",X"03",X"03",X"19",X"ec",X"4d",X"0b",X"4d",X"2e",X"2e",X"75",X"1b",X"0b",X"1b",X"3c",X"3c",X"0b",X"3c",X"0b",X"3c",X"1b",X"0b",X"0b",X"75",X"2e",X"2e",X"4d",X"1b",X"75",X"2e",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"71",X"19",X"03",X"19",X"71",X"2e",X"3c",X"1b",X"2e",X"03",X"21",X"1b",X"00",X"2e",X"ec",X"2e",X"1b",X"00",X"2e",X"2e",X"ec",X"14",X"2e",X"2e",X"03",X"03",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"2e",X"2e",X"fb",X"f4",X"fb",X"2e",X"2e",X"2e",X"fb",X"f4",X"00",X"00",X"2e",X"fb",X"00",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"92",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"1a",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"71",X"19",X"03",X"75",X"03",X"19",X"03",X"b2",X"27",X"75",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"03",X"75",X"03",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"d8",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"71",X"19",X"03",X"19",X"71",X"03",X"19",X"03",X"b2",X"03",X"75",X"03",X"19",X"03",X"1a",X"03",X"0b",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"7c",X"aa",X"61",X"0b",X"0b",X"1b",X"61",X"03",X"19",X"71",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"19",X"b2",X"19",X"3c",X"3c",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"2e",X"4d",X"1b",X"75",X"2e",X"ec",X"19",X"0b",X"3c",X"1a",X"1a",X"1a",X"3c",X"1b",X"75",X"03",X"1a",X"1b",X"1b",X"75",X"2e",X"ec",X"e9",X"3c",X"75",X"2e",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"ec",X"0b",X"0b",X"2e",X"19",X"2e",X"0b",X"0b",X"2e",X"2e",X"2e",X"0b",X"0b",X"2e",X"09",X"09",X"14",X"2e",X"1b",X"2e",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"03",X"1a",X"03",X"b2",X"19",X"71",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"fb",X"00",X"2e",X"fb",X"f4",X"3c",X"00",X"00",X"2e",X"fb",X"00",X"00",X"00",X"f4",X"00",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",X"60",X"aa",X"42",X"9e",X"98",X"0b",X"1b",X"0b",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"71",X"03",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"75",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"b2",X"27",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"19",X"71",X"19",X"03",X"1a",X"03",X"71",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"03",X"1a",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"9e",X"aa",X"60",X"98",X"0b",X"1b",X"0b",X"2f",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"0b",X"0b",X"0b",X"03",X"b2",X"03",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"30",X"e9",X"3c",X"19",X"2e",X"2e",X"4d",X"1b",X"1b",X"51",X"62",X"62",X"5d",X"0b",X"f5",X"3d",X"cf",X"3d",X"1b",X"00",X"2e",X"2e",X"25",X"00",X"3c",X"2e",X"2e",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"75",X"03",X"b2",X"03",X"2e",X"0b",X"1b",X"ec",X"03",X"2e",X"3c",X"0b",X"ec",X"2e",X"2e",X"1b",X"3c",X"2e",X"09",X"14",X"03",X"2e",X"0b",X"3c",X"2e",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"19",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"2e",X"f4",X"3c",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"3c",X"00",X"00",X"fb",X"00",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"aa",X"2c",X"aa",X"98",X"1b",X"0b",X"0b",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"71",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"71",X"19",X"03",X"75",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"19",X"03",X"19",X"71",X"19",X"71",X"03",X"03",X"1a",X"03",X"71",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"19",X"0b",X"0b",X"1b",X"17",X"6d",X"3f",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"79",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"75",X"03",X"1a",X"03",X"3c",X"2e",X"3c",X"19",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"03",X"19",X"b2",X"27",X"2e",X"25",X"00",X"0b",X"2e",X"2e",X"4d",X"0b",X"00",X"62",X"62",X"62",X"62",X"5d",X"cf",X"3d",X"25",X"3d",X"5d",X"0b",X"2e",X"ec",X"2e",X"1b",X"0b",X"3c",X"ea",X"2e",X"03",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"ec",X"0b",X"00",X"25",X"ec",X"2e",X"1b",X"0b",X"2e",X"2e",X"2e",X"3c",X"0b",X"2e",X"09",X"14",X"d8",X"2e",X"3c",X"0b",X"2e",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"19",X"71",X"19",X"b2",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"2e",X"fb",X"f4",X"91",X"f4",X"2e",X"2e",X"2e",X"fb",X"f4",X"00",X"00",X"fb",X"f4",X"00",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"79",X"6d",X"3f",X"6d",X"aa",X"12",X"aa",X"12",X"98",X"0b",X"0b",X"1b",X"d8",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"19",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"71",X"19",X"03",X"75",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"75",X"03",X"1a",X"03",X"75",X"03",X"1a",X"03",X"b2",X"27",X"1a",X"03",X"03",X"19",X"b2",X"27",X"19",X"03",X"03",X"b2",X"27",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"9e",X"aa",X"33",X"0b",X"0b",X"0b",X"2f",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"0b",X"2e",X"3c",X"1b",X"3c",X"0b",X"1b",X"0b",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"e5",X"1b",X"0b",X"3c",X"2e",X"ec",X"3d",X"5d",X"0b",X"51",X"15",X"cf",X"62",X"62",X"3d",X"3d",X"cf",X"3d",X"3a",X"1b",X"2e",X"2e",X"2e",X"1a",X"3c",X"1b",X"0b",X"00",X"2e",X"19",X"71",X"19",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"2e",X"1b",X"0b",X"25",X"ec",X"2e",X"3c",X"0b",X"2e",X"2e",X"ec",X"0b",X"1b",X"2e",X"14",X"03",X"03",X"2e",X"1b",X"0b",X"2e",X"03",X"19",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"fb",X"2e",X"fb",X"f4",X"fb",X"00",X"00",X"00",X"2e",X"fb",X"00",X"f4",X"fb",X"f4",X"fb",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"3b",X"6d",X"f0",X"6d",X"f0",X"60",X"aa",X"2c",X"aa",X"98",X"0b",X"1b",X"0b",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"03",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"75",X"03",X"b2",X"27",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"1a",X"03",X"03",X"75",X"03",X"75",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"27",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"19",X"0b",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"7c",X"61",X"0b",X"1b",X"83",X"2f",X"19",X"03",X"1a",X"03",X"03",X"19",X"71",X"19",X"03",X"03",X"03",X"19",X"03",X"1a",X"03",X"1b",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"00",X"03",X"b2",X"03",X"19",X"03",X"1a",X"2e",X"00",X"0b",X"3c",X"0b",X"2e",X"2e",X"e9",X"1b",X"0b",X"62",X"62",X"62",X"cf",X"3d",X"cf",X"f5",X"3d",X"3d",X"3d",X"5d",X"2e",X"ec",X"2e",X"51",X"75",X"e4",X"0b",X"0b",X"0b",X"2e",X"03",X"19",X"71",X"27",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"71",X"19",X"03",X"1a",X"03",X"b2",X"2e",X"0b",X"3c",X"4d",X"2e",X"2e",X"1b",X"3c",X"30",X"2e",X"2e",X"75",X"3c",X"2e",X"d8",X"03",X"03",X"2e",X"0b",X"3c",X"2e",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"71",X"19",X"71",X"19",X"71",X"19",X"03",X"03",X"1a",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f4",X"fb",X"2e",X"fb",X"f4",X"fb",X"f4",X"4f",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"f4",X"3c",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"aa",X"12",X"aa",X"98",X"0b",X"0b",X"0b",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"03",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"1b",X"0b",X"0b",X"53",X"54",X"3f",X"6d",X"3f",
    X"aa",X"9e",X"aa",X"9e",X"98",X"0b",X"0b",X"1b",X"ed",X"03",X"b2",X"27",X"19",X"b2",X"27",X"75",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"3c",X"2e",X"1b",X"0b",X"00",X"1b",X"0b",X"0b",X"03",X"1a",X"03",X"b2",X"03",X"2e",X"3c",X"0b",X"0b",X"0b",X"00",X"2e",X"2e",X"ec",X"0b",X"3c",X"62",X"51",X"62",X"62",X"62",X"3d",X"f5",X"3d",X"3d",X"3d",X"3d",X"ec",X"2e",X"2e",X"e9",X"3d",X"cf",X"3c",X"1b",X"0b",X"3c",X"2e",X"2e",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"cc",X"3c",X"1b",X"4d",X"2e",X"2e",X"3c",X"0b",X"e9",X"30",X"2e",X"19",X"0b",X"3d",X"2e",X"03",X"03",X"21",X"3c",X"0b",X"2e",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"b2",X"27",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"27",X"1a",X"03",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f4",X"fb",X"f4",X"2e",X"fb",X"f4",X"fb",X"f4",X"fb",X"fb",X"f4",X"fb",X"2e",X"fb",X"f4",X"91",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"7c",X"9e",X"aa",X"84",X"0b",X"0b",X"1b",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"75",X"03",X"b2",X"03",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"19",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"19",X"71",X"27",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"03",X"b2",X"27",X"19",X"03",X"0b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"2f",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"0b",X"2e",X"0b",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"03",X"2e",X"1b",X"0b",X"1b",X"15",X"3c",X"0b",X"2e",X"2e",X"2e",X"1b",X"0b",X"62",X"62",X"62",X"62",X"cf",X"3d",X"cf",X"25",X"cf",X"3d",X"3d",X"3d",X"30",X"ec",X"3d",X"3d",X"3d",X"e9",X"5d",X"3c",X"1b",X"0b",X"19",X"2e",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"71",X"19",X"b2",X"27",X"19",X"03",X"b2",X"03",X"2e",X"19",X"0b",X"75",X"2e",X"2e",X"3c",X"0b",X"3d",X"2e",X"ec",X"75",X"1b",X"25",X"ec",X"03",X"03",X"2e",X"0b",X"3c",X"2e",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"fb",X"f4",X"fb",X"f4",X"2e",X"2e",X"fb",X"f4",X"fb",X"f4",X"2e",X"2e",X"fb",X"f4",X"fb",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",X"60",X"aa",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"b2",X"27",X"19",X"71",X"75",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"b2",X"27",X"19",X"1a",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"75",X"03",X"03",X"1a",X"03",X"75",X"03",X"03",X"b2",X"19",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"19",X"3c",X"0b",X"3c",X"33",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"7c",X"9e",X"98",X"1b",X"0b",X"1b",X"61",X"03",X"b2",X"27",X"03",X"1a",X"03",X"03",X"75",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"3c",X"0b",X"3c",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"ec",X"0b",X"00",X"3a",X"51",X"3c",X"1b",X"51",X"ec",X"2e",X"0b",X"00",X"51",X"62",X"cf",X"3d",X"f5",X"f5",X"3d",X"cf",X"e9",X"3d",X"3d",X"3d",X"3d",X"ec",X"3d",X"3d",X"e9",X"3d",X"3d",X"5d",X"1b",X"3c",X"0b",X"1a",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"71",X"19",X"71",X"19",X"03",X"2e",X"75",X"0b",X"75",X"2e",X"3c",X"0b",X"0b",X"4d",X"2e",X"2e",X"19",X"0b",X"4d",X"2e",X"03",X"b2",X"2e",X"1b",X"0b",X"2e",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"2e",X"2e",X"2e",X"2e",X"fb",X"f4",X"fb",X"fb",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"60",X"aa",X"7c",X"33",X"0b",X"0b",X"0b",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"75",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"27",X"19",X"03",X"2e",X"ec",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"2e",X"2e",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"b2",X"19",X"71",X"27",X"19",X"1a",X"03",X"03",X"03",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"71",X"03",X"1a",X"03",X"0b",X"0b",X"0b",X"98",X"6d",X"3f",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"0b",X"0b",X"2f",X"03",X"19",X"71",X"19",X"03",X"b2",X"19",X"71",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"2e",X"0b",X"1b",X"0b",X"51",X"15",X"51",X"3c",X"51",X"15",X"30",X"1b",X"0b",X"62",X"62",X"15",X"cf",X"f5",X"3d",X"cf",X"25",X"cf",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"62",X"5d",X"1b",X"0b",X"3c",X"2e",X"19",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"2e",X"19",X"3c",X"75",X"0b",X"0b",X"3c",X"1b",X"4d",X"2e",X"2e",X"75",X"3c",X"4d",X"2e",X"03",X"19",X"2e",X"00",X"0b",X"2e",X"03",X"e5",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"f4",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"fb",X"f4",X"fb",X"f4",X"f4",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"aa",X"9e",X"98",X"1b",X"0b",X"1b",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"06",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"71",X"75",X"03",X"03",X"1a",X"03",X"b2",X"03",X"21",X"03",X"75",X"19",X"28",X"f0",X"f0",X"79",X"61",X"77",X"79",X"79",X"79",X"79",X"61",X"79",X"f0",X"98",X"2f",X"f0",X"98",X"79",X"f0",X"f0",X"75",X"19",X"03",X"21",X"2e",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"71",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"0b",X"1b",X"0b",X"3b",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"60",X"98",X"1b",X"0b",X"1b",X"79",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"d8",X"19",X"71",X"19",X"03",X"1a",X"03",X"19",X"2e",X"3c",X"3c",X"51",X"15",X"3a",X"51",X"15",X"3a",X"51",X"51",X"00",X"1b",X"51",X"62",X"62",X"62",X"3d",X"cf",X"f5",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"3d",X"5d",X"3c",X"1b",X"0b",X"2e",X"03",X"1a",X"03",X"03",X"b2",X"03",X"75",X"03",X"03",X"b2",X"03",X"19",X"ec",X"4d",X"0b",X"1b",X"0b",X"3c",X"0b",X"0b",X"75",X"2e",X"ec",X"19",X"0b",X"75",X"3c",X"2e",X"ec",X"2e",X"0b",X"00",X"4d",X"2e",X"1b",X"2e",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"d8",X"75",X"03",X"b2",X"03",X"19",X"03",X"b2",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"12",X"aa",X"7c",X"61",X"0b",X"0b",X"0b",X"75",X"03",X"b2",X"03",X"b2",X"03",X"03",X"03",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"cc",X"19",X"19",X"75",X"62",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"cf",X"15",X"62",X"cf",X"15",X"62",X"cf",X"15",X"51",X"f5",X"15",X"19",X"03",X"21",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"19",X"03",X"19",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"0b",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"9e",X"aa",X"84",X"0b",X"0b",X"0b",X"2f",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"27",X"19",X"03",X"b2",X"03",X"03",X"b2",X"2e",X"0b",X"0b",X"51",X"3a",X"15",X"51",X"51",X"15",X"51",X"15",X"0b",X"0b",X"62",X"62",X"62",X"62",X"cf",X"3d",X"3d",X"3d",X"cf",X"25",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"5d",X"1b",X"0b",X"1b",X"2e",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"d8",X"1a",X"03",X"b2",X"2e",X"4d",X"1b",X"3c",X"42",X"1a",X"e4",X"3c",X"75",X"2e",X"2e",X"4d",X"1b",X"75",X"0b",X"0b",X"0b",X"2e",X"1b",X"0b",X"00",X"3c",X"0b",X"30",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"91",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"3b",X"6d",X"3f",X"6d",X"f0",X"2c",X"aa",X"12",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"03",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"75",X"03",X"2e",X"03",X"28",X"62",X"51",X"62",X"15",X"cf",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"15",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"15",X"51",X"f5",X"75",X"19",X"2e",X"03",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"71",X"03",X"03",X"b2",X"03",X"75",X"03",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"7c",X"61",X"0b",X"1b",X"0b",X"79",X"03",X"b2",X"03",X"1a",X"03",X"03",X"75",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"21",X"1b",X"1b",X"3a",X"15",X"51",X"51",X"15",X"3a",X"51",X"15",X"51",X"3c",X"1b",X"51",X"62",X"cf",X"62",X"3d",X"f5",X"cf",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"e9",X"3d",X"5d",X"3c",X"0b",X"1b",X"2e",X"03",X"19",X"71",X"03",X"03",X"19",X"b2",X"27",X"19",X"03",X"30",X"e9",X"00",X"0b",X"ea",X"ea",X"1a",X"1b",X"75",X"2e",X"2e",X"4d",X"1b",X"75",X"3c",X"0b",X"1b",X"0b",X"3c",X"0b",X"0b",X"0b",X"0b",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"aa",X"2c",X"aa",X"ba",X"0b",X"0b",X"1b",X"1a",X"03",X"b2",X"27",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"03",X"21",X"75",X"62",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"15",X"62",X"75",X"ec",X"27",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"75",X"03",X"1a",X"03",X"03",X"b2",X"ad",X"1b",X"0b",X"53",X"6d",X"3f",X"6d",X"f0",
    X"9e",X"aa",X"9e",X"aa",X"98",X"0b",X"0b",X"0b",X"2f",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"19",X"71",X"03",X"1a",X"03",X"75",X"03",X"03",X"b2",X"03",X"19",X"2e",X"0b",X"3c",X"51",X"51",X"15",X"3a",X"51",X"15",X"51",X"3a",X"62",X"3c",X"0b",X"62",X"62",X"15",X"cf",X"62",X"cf",X"25",X"3d",X"cf",X"e9",X"3d",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"e9",X"3d",X"3d",X"3d",X"e9",X"3d",X"5d",X"1b",X"3c",X"0b",X"2e",X"2e",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"2e",X"25",X"1b",X"3c",X"ea",X"19",X"1a",X"3c",X"1a",X"ec",X"2e",X"e9",X"00",X"19",X"0b",X"1b",X"0b",X"00",X"0b",X"0b",X"3c",X"0b",X"3c",X"2e",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"4a",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"79",X"6d",X"f0",X"6d",X"aa",X"12",X"aa",X"9e",X"98",X"0b",X"1b",X"0b",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"75",X"03",X"b2",X"03",X"1a",X"03",X"03",X"19",X"b2",X"19",X"03",X"2e",X"19",X"15",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"cf",X"15",X"62",X"51",X"62",X"62",X"cf",X"15",X"51",X"62",X"15",X"f5",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"19",X"ec",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"19",X"3c",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"aa",X"7c",X"aa",X"84",X"0b",X"1b",X"0b",X"79",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"03",X"75",X"03",X"b2",X"03",X"03",X"b2",X"27",X"03",X"1a",X"03",X"03",X"71",X"19",X"71",X"19",X"03",X"2e",X"0b",X"00",X"0b",X"3a",X"15",X"51",X"15",X"3a",X"51",X"51",X"15",X"51",X"00",X"3c",X"51",X"62",X"f5",X"62",X"f5",X"3d",X"cf",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"e9",X"3d",X"5d",X"3c",X"0b",X"00",X"ea",X"2e",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"ec",X"0b",X"0b",X"19",X"42",X"75",X"0b",X"0b",X"2e",X"ec",X"25",X"1b",X"1a",X"75",X"b2",X"0b",X"1b",X"0b",X"00",X"0b",X"3c",X"0b",X"2e",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"19",X"00",X"00",X"f4",X"3c",X"8f",X"4f",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"53",X"6d",X"f0",X"6d",X"3f",X"2c",X"aa",X"7c",X"aa",X"98",X"0b",X"0b",X"0b",X"19",X"71",X"19",X"03",X"19",X"71",X"19",X"b2",X"03",X"03",X"03",X"1a",X"03",X"03",X"75",X"03",X"b2",X"27",X"19",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"75",X"03",X"19",X"71",X"19",X"b2",X"03",X"03",X"b2",X"2e",X"1a",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"cf",X"62",X"51",X"62",X"15",X"f5",X"62",X"62",X"cf",X"15",X"62",X"62",X"cf",X"15",X"62",X"51",X"62",X"62",X"62",X"51",X"1a",X"2e",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"75",X"03",X"03",X"b2",X"03",X"03",X"19",X"03",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"19",X"1a",X"03",X"03",X"0b",X"0b",X"0b",X"3b",X"6d",X"f0",X"6d",X"3f",
    X"60",X"aa",X"12",X"aa",X"98",X"83",X"0b",X"0b",X"2f",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"2e",X"1b",X"0b",X"15",X"51",X"51",X"51",X"51",X"15",X"3a",X"15",X"51",X"15",X"51",X"1b",X"62",X"62",X"15",X"cf",X"3d",X"f5",X"cf",X"25",X"cf",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"5d",X"1b",X"0b",X"00",X"1a",X"2e",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"2e",X"3c",X"0b",X"ea",X"ea",X"ea",X"3c",X"1b",X"2e",X"2e",X"2e",X"3c",X"b2",X"19",X"75",X"19",X"b2",X"0b",X"1b",X"0b",X"0b",X"00",X"2e",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"f4",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"9e",X"aa",X"9e",X"98",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"b2",X"27",X"75",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"27",X"19",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"2e",X"2f",X"62",X"62",X"15",X"f5",X"15",X"f5",X"cf",X"15",X"62",X"51",X"62",X"62",X"15",X"f5",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"cf",X"62",X"15",X"cf",X"15",X"62",X"79",X"2e",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"d8",X"75",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"1b",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"aa",X"2c",X"aa",X"33",X"1b",X"0b",X"0b",X"79",X"03",X"71",X"19",X"b2",X"03",X"1a",X"03",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"ec",X"0b",X"3c",X"51",X"15",X"3a",X"15",X"51",X"51",X"51",X"51",X"51",X"51",X"15",X"cf",X"62",X"51",X"62",X"62",X"62",X"cf",X"f5",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"3d",X"3d",X"e9",X"3d",X"3d",X"3d",X"e9",X"3d",X"3d",X"e9",X"15",X"3c",X"0b",X"0b",X"3c",X"2e",X"03",X"75",X"03",X"03",X"19",X"71",X"2e",X"0b",X"3c",X"ea",X"ea",X"75",X"0b",X"0b",X"2e",X"2e",X"2e",X"1b",X"1a",X"75",X"75",X"19",X"1a",X"0b",X"00",X"0b",X"3c",X"0b",X"2e",X"03",X"19",X"03",X"b2",X"27",X"75",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"19",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"9e",X"aa",X"7c",X"aa",X"74",X"0b",X"0b",X"1b",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"71",X"19",X"03",X"19",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"2e",X"2f",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"15",X"62",X"51",X"62",X"15",X"f5",X"62",X"15",X"62",X"62",X"62",X"51",X"62",X"15",X"51",X"62",X"62",X"15",X"f5",X"51",X"62",X"62",X"77",X"2e",X"03",X"75",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"75",X"03",X"03",X"1a",X"03",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"12",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"2f",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"19",X"71",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"19",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"2e",X"0b",X"0b",X"3a",X"51",X"15",X"3a",X"51",X"15",X"3a",X"15",X"51",X"15",X"51",X"62",X"62",X"15",X"62",X"cf",X"3d",X"f5",X"3d",X"3d",X"cf",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"e9",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"e9",X"4d",X"5d",X"3c",X"0b",X"0b",X"2e",X"2e",X"03",X"1a",X"71",X"19",X"2e",X"3c",X"0b",X"ea",X"ea",X"ea",X"3c",X"1b",X"2e",X"ec",X"2e",X"3c",X"0b",X"19",X"75",X"19",X"75",X"1b",X"0b",X"0b",X"0b",X"3c",X"2e",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"00",X"00",X"fb",X"00",X"a4",X"91",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"3b",X"6d",X"3f",X"f0",X"6d",X"aa",X"aa",X"60",X"aa",X"98",X"0b",X"0b",X"1b",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"2e",X"98",X"62",X"62",X"15",X"62",X"62",X"15",X"62",X"51",X"62",X"cf",X"62",X"62",X"62",X"cf",X"15",X"51",X"cf",X"62",X"51",X"15",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"79",X"2e",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"71",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"71",X"03",X"b2",X"19",X"03",X"b2",X"83",X"3c",X"0b",X"53",X"6d",X"f0",X"6d",X"3f",
    X"9e",X"aa",X"7c",X"9e",X"98",X"0b",X"1b",X"83",X"2f",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"03",X"75",X"03",X"03",X"b2",X"27",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"ec",X"0b",X"3c",X"15",X"51",X"51",X"51",X"15",X"51",X"51",X"51",X"51",X"15",X"62",X"51",X"f5",X"51",X"62",X"62",X"cf",X"3d",X"f5",X"cf",X"e9",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"5d",X"3c",X"0b",X"3c",X"ea",X"2e",X"03",X"19",X"03",X"21",X"1b",X"0b",X"19",X"ea",X"75",X"0b",X"0b",X"2e",X"2e",X"2e",X"3c",X"0b",X"75",X"75",X"19",X"75",X"0b",X"1b",X"0b",X"00",X"0b",X"2e",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"d8",X"19",X"71",X"19",X"b2",X"27",X"19",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f4",X"fb",X"f4",X"fb",X"91",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"4f",X"f4",X"fb",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"6d",X"aa",X"12",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"d8",X"19",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"75",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"ec",X"2f",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"62",X"62",X"cf",X"15",X"62",X"cf",X"15",X"f5",X"15",X"62",X"62",X"51",X"62",X"ed",X"2e",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"19",X"03",X"19",X"03",X"71",X"19",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"2c",X"aa",X"aa",X"98",X"0b",X"0b",X"0b",X"2f",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"19",X"71",X"27",X"1a",X"03",X"b2",X"27",X"19",X"71",X"19",X"71",X"19",X"71",X"19",X"03",X"03",X"e5",X"3c",X"0b",X"51",X"15",X"3a",X"15",X"3a",X"51",X"15",X"3a",X"15",X"51",X"51",X"15",X"62",X"15",X"62",X"62",X"62",X"3d",X"cf",X"3d",X"f5",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"e9",X"3d",X"e9",X"4d",X"4d",X"5d",X"3c",X"0b",X"1b",X"1a",X"2e",X"2e",X"03",X"2e",X"0b",X"00",X"42",X"19",X"42",X"1b",X"1b",X"75",X"2e",X"2e",X"3c",X"0b",X"75",X"19",X"75",X"75",X"3c",X"0b",X"3c",X"0b",X"0b",X"2e",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"b2",X"27",X"19",X"03",X"03",X"b2",X"03",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"f4",X"fb",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"2c",X"aa",X"12",X"98",X"0b",X"0b",X"0b",X"19",X"71",X"19",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"19",X"71",X"27",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"2e",X"54",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"51",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"cf",X"15",X"62",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"d8",X"75",X"03",X"19",X"03",X"19",X"03",X"b2",X"d8",X"19",X"71",X"19",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"0b",X"0b",X"0b",X"3b",X"f0",X"6d",X"3f",X"6d",
    X"aa",X"12",X"aa",X"9e",X"98",X"1b",X"0b",X"0b",X"79",X"03",X"19",X"03",X"b2",X"27",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"19",X"03",X"19",X"03",X"b2",X"2e",X"1b",X"0b",X"3a",X"51",X"51",X"51",X"15",X"51",X"51",X"15",X"51",X"51",X"15",X"f5",X"62",X"cf",X"62",X"62",X"62",X"cf",X"3d",X"f5",X"3d",X"cf",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"3d",X"e9",X"4d",X"3d",X"e9",X"4d",X"4d",X"bf",X"3c",X"3c",X"0b",X"0b",X"3c",X"2e",X"2e",X"1b",X"0b",X"ea",X"ea",X"75",X"ea",X"0b",X"75",X"19",X"2e",X"1b",X"0b",X"19",X"75",X"75",X"19",X"0b",X"0b",X"00",X"0b",X"1b",X"2e",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f4",X"4f",X"f4",X"4f",X"f4",X"fb",X"00",X"00",X"00",X"00",X"fb",X"f4",X"fb",X"91",X"f4",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",X"9e",X"aa",X"9e",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"75",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"19",X"03",X"2e",X"2f",X"62",X"51",X"62",X"51",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"cf",X"62",X"15",X"f5",X"51",X"62",X"62",X"15",X"62",X"62",X"62",X"51",X"62",X"51",X"79",X"2e",X"1a",X"03",X"19",X"03",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"d8",X"03",X"b2",X"03",X"b2",X"27",X"19",X"b2",X"27",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"19",X"3c",X"0b",X"00",X"98",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"6d",X"aa",X"7c",X"61",X"0b",X"0b",X"1b",X"2f",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"b2",X"19",X"b2",X"27",X"19",X"71",X"27",X"19",X"03",X"19",X"71",X"19",X"b2",X"03",X"b2",X"03",X"19",X"2e",X"3c",X"0b",X"15",X"51",X"15",X"3a",X"51",X"15",X"3a",X"51",X"51",X"15",X"51",X"15",X"51",X"62",X"51",X"cf",X"62",X"f5",X"3d",X"cf",X"25",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"3d",X"3d",X"3d",X"e9",X"4d",X"3d",X"e9",X"4d",X"4d",X"4d",X"e9",X"4d",X"5d",X"0b",X"3c",X"0b",X"0b",X"30",X"0b",X"1b",X"ea",X"19",X"ea",X"75",X"ea",X"19",X"1a",X"75",X"0b",X"1b",X"75",X"75",X"19",X"75",X"0b",X"1b",X"0b",X"0b",X"3c",X"2e",X"75",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"71",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f4",X"00",X"00",X"f4",X"00",X"00",X"fb",X"f4",X"91",X"f4",X"00",X"3c",X"f4",X"fb",X"f4",X"91",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"3f",X"f0",X"7c",X"aa",X"7c",X"aa",X"61",X"0b",X"0b",X"0b",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"71",X"27",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"e5",X"2f",X"62",X"15",X"f5",X"62",X"62",X"51",X"62",X"cf",X"15",X"62",X"62",X"cf",X"15",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"15",X"f5",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"ed",X"2e",X"03",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"19",X"03",X"b2",X"03",X"b2",X"1b",X"83",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"36",X"9e",X"aa",X"98",X"1b",X"83",X"0b",X"2f",X"19",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"b2",X"2e",X"1b",X"0b",X"0b",X"3a",X"51",X"15",X"51",X"51",X"51",X"15",X"51",X"51",X"62",X"62",X"62",X"15",X"f5",X"62",X"62",X"3d",X"cf",X"f5",X"3d",X"cf",X"25",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"e9",X"4d",X"3d",X"4d",X"4d",X"4d",X"5d",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"19",X"42",X"19",X"ea",X"75",X"75",X"19",X"19",X"b2",X"0b",X"75",X"19",X"75",X"19",X"b2",X"0b",X"3c",X"0b",X"00",X"2e",X"19",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"71",X"19",X"b2",X"03",X"03",X"03",X"b2",X"03",X"19",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"fb",X"2e",X"fb",X"00",X"fb",X"f4",X"3c",X"f4",X"fb",X"f4",X"fb",X"f4",X"00",X"fb",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"6d",X"6d",X"9e",X"aa",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"03",X"b2",X"27",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"75",X"03",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"b2",X"27",X"75",X"03",X"2e",X"98",X"62",X"62",X"51",X"15",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"cf",X"62",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"15",X"cf",X"62",X"15",X"62",X"62",X"15",X"62",X"51",X"f0",X"2e",X"03",X"1a",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"71",X"19",X"03",X"19",X"0b",X"1b",X"0b",X"3b",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"60",X"aa",X"60",X"98",X"0b",X"1b",X"0b",X"79",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"b2",X"19",X"03",X"03",X"1a",X"ec",X"0b",X"3c",X"51",X"15",X"3a",X"51",X"15",X"51",X"3a",X"15",X"51",X"15",X"51",X"62",X"cf",X"15",X"f5",X"62",X"cf",X"3d",X"3d",X"f5",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"e9",X"4d",X"4d",X"4d",X"e9",X"4d",X"4d",X"4d",X"1b",X"1b",X"0b",X"00",X"0b",X"0b",X"19",X"ea",X"ea",X"75",X"ea",X"19",X"75",X"75",X"1a",X"1b",X"75",X"19",X"75",X"75",X"1a",X"1b",X"0b",X"0b",X"1b",X"2e",X"4d",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f4",X"fb",X"2e",X"f4",X"00",X"fb",X"f4",X"00",X"fb",X"f4",X"91",X"f4",X"00",X"fb",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"f0",X"3f",X"f0",X"aa",X"aa",X"92",X"aa",X"98",X"0b",X"0b",X"1b",X"d8",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"b2",X"19",X"71",X"19",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"21",X"2f",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"51",X"62",X"51",X"cf",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"cf",X"62",X"51",X"62",X"62",X"2f",X"2e",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"aa",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"2f",X"03",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"19",X"03",X"71",X"19",X"03",X"2e",X"1b",X"0b",X"3a",X"51",X"15",X"3a",X"51",X"15",X"51",X"51",X"15",X"51",X"62",X"62",X"51",X"62",X"15",X"cf",X"3d",X"f5",X"cf",X"3d",X"15",X"3c",X"0b",X"0b",X"00",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"e9",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"3d",X"4d",X"1b",X"0b",X"0b",X"00",X"0b",X"19",X"42",X"75",X"ea",X"19",X"75",X"75",X"19",X"b2",X"0b",X"19",X"75",X"75",X"19",X"b2",X"0b",X"3c",X"0b",X"3c",X"3d",X"4d",X"03",X"1a",X"03",X"03",X"b2",X"03",X"75",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f4",X"fb",X"f4",X"fb",X"fb",X"f4",X"2e",X"00",X"fb",X"f4",X"fb",X"f4",X"fb",X"00",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"6d",X"aa",X"60",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"2e",X"54",X"62",X"62",X"15",X"cf",X"62",X"51",X"62",X"62",X"15",X"cf",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"62",X"51",X"15",X"62",X"62",X"51",X"62",X"62",X"15",X"f5",X"cf",X"15",X"98",X"2e",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"75",X"03",X"1a",X"03",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"0b",X"1b",X"0b",X"3b",X"1a",X"6d",X"f0",X"6d",
    X"9e",X"7c",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"79",X"03",X"b2",X"19",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"2e",X"00",X"0b",X"15",X"51",X"51",X"15",X"3a",X"51",X"15",X"51",X"51",X"15",X"51",X"62",X"62",X"62",X"62",X"62",X"62",X"cf",X"3d",X"51",X"3c",X"0b",X"1b",X"0b",X"0b",X"1b",X"3d",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"e9",X"3d",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"e9",X"4d",X"4d",X"e9",X"4d",X"19",X"4d",X"1b",X"1b",X"0b",X"00",X"42",X"19",X"ea",X"75",X"42",X"75",X"19",X"75",X"1a",X"e4",X"b2",X"19",X"75",X"19",X"1a",X"00",X"0b",X"0b",X"00",X"25",X"4d",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f4",X"4f",X"2e",X"fb",X"f4",X"2e",X"2e",X"fb",X"f4",X"fb",X"f4",X"91",X"f4",X"00",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"3f",X"aa",X"9e",X"aa",X"60",X"61",X"0b",X"0b",X"0b",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"2e",X"2f",X"f5",X"51",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"15",X"f5",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"cf",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"ed",X"2e",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"27",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"0b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"2f",X"1a",X"03",X"03",X"03",X"19",X"03",X"03",X"1a",X"03",X"19",X"b2",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"75",X"03",X"2e",X"0b",X"1b",X"51",X"15",X"3a",X"51",X"15",X"51",X"51",X"3a",X"15",X"51",X"51",X"15",X"51",X"62",X"51",X"cf",X"62",X"3d",X"f5",X"1b",X"0b",X"1b",X"0b",X"00",X"0b",X"00",X"0b",X"3d",X"3d",X"3d",X"e9",X"3d",X"3d",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"e9",X"3d",X"e9",X"4d",X"4d",X"4d",X"4d",X"4d",X"19",X"4d",X"19",X"42",X"1a",X"e4",X"0b",X"19",X"ea",X"bf",X"19",X"75",X"19",X"75",X"19",X"06",X"0b",X"1a",X"75",X"19",X"75",X"b2",X"0b",X"1b",X"0b",X"0b",X"4d",X"e9",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"19",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"fb",X"f4",X"2e",X"2e",X"2e",X"2e",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"00",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"3b",X"6d",X"f0",X"6d",X"6d",X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"0b",X"3c",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"19",X"b2",X"27",X"19",X"03",X"b2",X"2e",X"2f",X"62",X"62",X"15",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"f5",X"15",X"cf",X"15",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"62",X"cf",X"62",X"62",X"62",X"15",X"62",X"51",X"61",X"2e",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"0b",X"0b",X"1b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"12",X"98",X"0b",X"0b",X"1b",X"61",X"03",X"03",X"b2",X"19",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"75",X"03",X"b2",X"27",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"2e",X"3c",X"0b",X"3a",X"51",X"15",X"3a",X"51",X"51",X"15",X"51",X"51",X"15",X"62",X"62",X"62",X"15",X"62",X"51",X"3d",X"f5",X"cf",X"1b",X"0b",X"00",X"0b",X"2e",X"1b",X"0b",X"0b",X"3c",X"25",X"e9",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"e9",X"4d",X"3d",X"e9",X"4d",X"3d",X"4d",X"e9",X"4d",X"4d",X"4d",X"bf",X"ea",X"1a",X"1b",X"ea",X"ea",X"ea",X"19",X"ea",X"75",X"75",X"75",X"19",X"3c",X"b2",X"19",X"75",X"75",X"aa",X"1b",X"3c",X"0b",X"1b",X"4d",X"3d",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f4",X"fb",X"2e",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"91",X"f4",X"fb",X"f4",X"91",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"9e",X"aa",X"9e",X"98",X"1b",X"0b",X"0b",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"d8",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"2e",X"2f",X"62",X"51",X"62",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"62",X"cf",X"15",X"f5",X"62",X"62",X"cf",X"15",X"62",X"51",X"62",X"62",X"51",X"15",X"62",X"51",X"15",X"62",X"51",X"62",X"62",X"2f",X"2e",X"03",X"19",X"b2",X"27",X"19",X"03",X"1a",X"03",X"03",X"b2",X"d8",X"03",X"1a",X"71",X"19",X"03",X"1a",X"03",X"b2",X"27",X"1a",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"27",X"b2",X"03",X"19",X"03",X"0b",X"1b",X"0b",X"33",X"6d",X"3f",X"6d",X"f0",
    X"9e",X"aa",X"9e",X"aa",X"98",X"0b",X"1b",X"0b",X"2f",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"75",X"2e",X"3c",X"0b",X"15",X"51",X"15",X"51",X"15",X"3a",X"51",X"15",X"51",X"51",X"15",X"cf",X"62",X"62",X"62",X"62",X"cf",X"3d",X"f5",X"1b",X"0b",X"0b",X"3c",X"2e",X"1b",X"0b",X"3c",X"0b",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"e9",X"4d",X"4d",X"4d",X"e9",X"3d",X"4d",X"4d",X"4d",X"4d",X"ea",X"ea",X"ea",X"ea",X"ea",X"75",X"ea",X"75",X"19",X"75",X"19",X"75",X"0b",X"1a",X"19",X"75",X"19",X"75",X"3c",X"0b",X"0b",X"3c",X"75",X"2e",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f4",X"91",X"f4",X"2e",X"fb",X"f4",X"91",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"7c",X"aa",X"7c",X"61",X"0b",X"0b",X"1b",X"03",X"1a",X"03",X"19",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"2e",X"2f",X"62",X"62",X"51",X"62",X"51",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"cf",X"62",X"62",X"51",X"79",X"2e",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"b2",X"19",X"03",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"3f",
    X"aa",X"7c",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"79",X"03",X"19",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"27",X"2e",X"3c",X"0b",X"3a",X"51",X"3a",X"51",X"51",X"15",X"51",X"51",X"51",X"15",X"f5",X"51",X"62",X"cf",X"62",X"62",X"3d",X"cf",X"3d",X"0b",X"1b",X"0b",X"3c",X"2e",X"2e",X"3c",X"0b",X"1b",X"0b",X"3d",X"e9",X"e9",X"3d",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"e9",X"4d",X"4d",X"4d",X"4d",X"4d",X"3d",X"4d",X"fc",X"bf",X"ea",X"ea",X"ea",X"ea",X"ea",X"19",X"ea",X"75",X"19",X"75",X"aa",X"1b",X"b2",X"19",X"75",X"75",X"19",X"0b",X"0b",X"00",X"0b",X"75",X"2e",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"b2",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f4",X"fb",X"f4",X"2e",X"fb",X"f4",X"fb",X"f4",X"fb",X"fb",X"f4",X"fb",X"2e",X"fb",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"12",X"aa",X"aa",X"9e",X"54",X"1b",X"0b",X"1b",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"71",X"2e",X"98",X"51",X"62",X"62",X"62",X"15",X"f5",X"51",X"62",X"62",X"51",X"62",X"15",X"f5",X"62",X"51",X"1d",X"62",X"62",X"51",X"cf",X"15",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"15",X"62",X"62",X"54",X"2e",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"1b",X"0b",X"1b",X"17",X"6d",X"f0",X"6d",X"6d",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"2f",X"03",X"b2",X"03",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"03",X"21",X"1b",X"0b",X"51",X"15",X"15",X"3a",X"15",X"51",X"3a",X"15",X"62",X"51",X"15",X"62",X"51",X"15",X"62",X"62",X"cf",X"3d",X"3d",X"5d",X"0b",X"3c",X"0b",X"b2",X"2e",X"2e",X"ea",X"1b",X"0b",X"3c",X"25",X"3d",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"e9",X"4d",X"4d",X"4d",X"4d",X"e9",X"4d",X"4d",X"19",X"4d",X"fc",X"bf",X"ea",X"ea",X"ea",X"bf",X"ea",X"75",X"19",X"75",X"75",X"19",X"3c",X"1a",X"aa",X"75",X"19",X"1a",X"3c",X"1b",X"0b",X"0b",X"19",X"2e",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f4",X"fb",X"fb",X"f4",X"2e",X"2e",X"fb",X"f4",X"fb",X"f4",X"2e",X"2e",X"fb",X"f4",X"fb",X"f4",X"3c",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"3f",X"6d",X"aa",X"7c",X"aa",X"74",X"0b",X"0b",X"0b",X"03",X"03",X"1a",X"03",X"19",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"27",X"75",X"03",X"b2",X"27",X"19",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"d8",X"19",X"2e",X"2f",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"cf",X"15",X"f5",X"51",X"62",X"3a",X"18",X"8e",X"51",X"51",X"62",X"62",X"62",X"cf",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"ed",X"2e",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"71",X"19",X"71",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"f0",
    X"aa",X"7c",X"0d",X"60",X"61",X"0b",X"0b",X"83",X"2f",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"71",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"b2",X"19",X"2e",X"3c",X"3c",X"3a",X"51",X"51",X"3a",X"15",X"51",X"51",X"51",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"f5",X"cf",X"62",X"1b",X"0b",X"3c",X"1a",X"2e",X"03",X"cc",X"4d",X"0b",X"0b",X"3c",X"25",X"e9",X"3d",X"3d",X"e9",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"e9",X"4d",X"4d",X"4d",X"3d",X"4d",X"4d",X"ea",X"ea",X"ea",X"ea",X"42",X"19",X"ea",X"75",X"ea",X"19",X"75",X"19",X"75",X"0b",X"1b",X"75",X"19",X"75",X"19",X"0b",X"0b",X"00",X"0b",X"75",X"2e",X"03",X"b2",X"27",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"d8",X"03",X"19",X"03",X"b2",X"19",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"2e",X"2e",X"2e",X"2e",X"fb",X"f4",X"fb",X"f4",X"91",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"c6",X"6d",X"f0",X"6d",X"6d",X"aa",X"aa",X"9e",X"aa",X"98",X"1b",X"0b",X"1b",X"d8",X"1a",X"03",X"b2",X"27",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"2e",X"2f",X"62",X"51",X"15",X"cf",X"62",X"62",X"62",X"51",X"62",X"62",X"15",X"f5",X"51",X"8f",X"8e",X"8e",X"41",X"51",X"51",X"62",X"15",X"51",X"62",X"cf",X"62",X"15",X"51",X"62",X"51",X"62",X"62",X"61",X"2e",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"71",X"03",X"1a",X"03",X"19",X"03",X"75",X"03",X"1a",X"03",X"1a",X"03",X"03",X"19",X"00",X"0b",X"1b",X"3b",X"3f",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"7c",X"aa",X"98",X"0b",X"1b",X"0b",X"2f",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"e5",X"1b",X"0b",X"51",X"15",X"3a",X"15",X"51",X"15",X"51",X"15",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"cf",X"3d",X"3d",X"3d",X"1b",X"0b",X"0b",X"0b",X"06",X"2e",X"03",X"21",X"2e",X"3c",X"0b",X"0b",X"3d",X"e9",X"e9",X"3d",X"3d",X"e9",X"3d",X"e9",X"4d",X"4d",X"4d",X"4d",X"4d",X"e9",X"4d",X"4d",X"bf",X"4d",X"ea",X"ea",X"ea",X"ea",X"ea",X"19",X"ea",X"75",X"75",X"19",X"75",X"75",X"0b",X"3c",X"1a",X"19",X"75",X"aa",X"3c",X"0b",X"00",X"0b",X"00",X"2e",X"03",X"19",X"b2",X"19",X"03",X"b2",X"03",X"b2",X"19",X"03",X"19",X"b2",X"19",X"b2",X"03",X"19",X"03",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"91",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"9e",X"7c",X"aa",X"60",X"98",X"0b",X"0b",X"0b",X"19",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"1a",X"2e",X"2f",X"62",X"62",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"18",X"8e",X"8e",X"8e",X"8e",X"8e",X"51",X"51",X"62",X"62",X"15",X"f5",X"51",X"62",X"62",X"62",X"15",X"51",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"83",X"0b",X"0b",X"98",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"9e",X"98",X"1b",X"0b",X"0b",X"79",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"19",X"71",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"03",X"19",X"b2",X"03",X"2e",X"ec",X"0b",X"1b",X"51",X"15",X"51",X"51",X"3a",X"51",X"15",X"62",X"51",X"cf",X"15",X"62",X"62",X"62",X"62",X"3d",X"cf",X"25",X"cf",X"e4",X"0b",X"3c",X"0b",X"2e",X"03",X"1a",X"03",X"2e",X"1b",X"0b",X"3c",X"25",X"3d",X"3d",X"e9",X"3d",X"e9",X"3d",X"e9",X"3d",X"4d",X"e9",X"4d",X"4d",X"4d",X"4d",X"4d",X"fc",X"bf",X"ea",X"ea",X"ea",X"ea",X"ea",X"75",X"ea",X"19",X"75",X"75",X"19",X"3c",X"0b",X"19",X"75",X"75",X"19",X"1b",X"0b",X"0b",X"1b",X"0b",X"2e",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"03",X"19",X"b2",X"03",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f4",X"91",X"f4",X"fb",X"f4",X"fb",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"91",X"f4",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"b2",X"27",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"2e",X"ed",X"62",X"62",X"51",X"62",X"62",X"cf",X"15",X"62",X"51",X"62",X"51",X"de",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"51",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"ed",X"2e",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"75",X"03",X"71",X"19",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"75",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"19",X"1b",X"0b",X"0b",X"3b",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"33",X"0b",X"0b",X"1b",X"2f",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"06",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"4d",X"3c",X"0b",X"51",X"3a",X"51",X"15",X"51",X"15",X"51",X"51",X"15",X"62",X"62",X"cf",X"15",X"62",X"62",X"cf",X"f5",X"3d",X"3d",X"5d",X"3c",X"0b",X"0b",X"3c",X"2e",X"03",X"1a",X"03",X"2e",X"3c",X"0b",X"0b",X"3a",X"e9",X"3d",X"3d",X"e9",X"3d",X"e9",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"bf",X"4d",X"fc",X"bf",X"ea",X"ea",X"ea",X"bf",X"19",X"19",X"75",X"75",X"19",X"75",X"0b",X"1b",X"75",X"75",X"19",X"75",X"1b",X"0b",X"3c",X"0b",X"3c",X"2e",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"00",X"00",X"f4",X"3c",X"8f",X"4f",X"f4",X"fb",X"f4",X"f4",X"91",X"f4",X"f4",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"fb",X"f4",X"4f",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"53",X"6d",X"f0",X"3f",X"6d",X"aa",X"6d",X"36",X"60",X"61",X"0b",X"0b",X"0b",X"19",X"71",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"d8",X"19",X"03",X"1a",X"2e",X"2f",X"f5",X"51",X"62",X"15",X"51",X"62",X"51",X"62",X"62",X"a1",X"18",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"51",X"51",X"62",X"51",X"62",X"cf",X"62",X"15",X"f5",X"51",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"27",X"03",X"1a",X"03",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"75",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"83",X"3c",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"9e",X"aa",X"9e",X"7c",X"61",X"0b",X"1b",X"0b",X"2f",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"2e",X"3c",X"3c",X"51",X"15",X"3a",X"51",X"51",X"51",X"15",X"62",X"62",X"51",X"62",X"62",X"cf",X"3d",X"62",X"3d",X"3d",X"cf",X"62",X"1b",X"0b",X"3c",X"0b",X"3c",X"2e",X"03",X"1a",X"03",X"2e",X"1b",X"0b",X"00",X"0b",X"25",X"e9",X"3d",X"e9",X"3d",X"e9",X"4d",X"3d",X"e9",X"3d",X"4d",X"4d",X"4d",X"42",X"19",X"fc",X"bf",X"ea",X"ea",X"ea",X"aa",X"ea",X"75",X"19",X"75",X"75",X"0b",X"3c",X"75",X"19",X"75",X"75",X"0b",X"00",X"0b",X"3c",X"0b",X"2e",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"75",X"03",X"1a",X"03",X"03",X"19",X"71",X"19",X"03",X"1a",X"00",X"00",X"fb",X"00",X"a4",X"4f",X"f4",X"4f",X"fb",X"fb",X"fb",X"fb",X"fb",X"91",X"f4",X"4f",X"fb",X"f4",X"4f",X"f4",X"fb",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"12",X"aa",X"9e",X"aa",X"98",X"0b",X"1b",X"0b",X"d8",X"1a",X"03",X"03",X"71",X"19",X"03",X"03",X"71",X"19",X"71",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"71",X"19",X"71",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"e5",X"2f",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"f5",X"51",X"18",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"a1",X"62",X"62",X"62",X"15",X"62",X"cf",X"15",X"62",X"51",X"79",X"2e",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"19",X"1b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"0b",X"0b",X"79",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"71",X"27",X"4d",X"1b",X"0b",X"51",X"3a",X"15",X"51",X"15",X"3a",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"cf",X"3d",X"cf",X"3d",X"25",X"3d",X"5d",X"00",X"0b",X"1b",X"0b",X"0b",X"ec",X"03",X"1a",X"03",X"2e",X"3c",X"0b",X"0b",X"00",X"3d",X"4d",X"e9",X"4d",X"4d",X"4d",X"4d",X"4d",X"e9",X"4d",X"4d",X"19",X"4d",X"ea",X"ea",X"19",X"42",X"19",X"19",X"19",X"75",X"19",X"75",X"75",X"19",X"1b",X"0b",X"75",X"aa",X"19",X"75",X"1b",X"0b",X"0b",X"0b",X"3c",X"2e",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"71",X"19",X"71",X"19",X"03",X"1a",X"03",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"7c",X"aa",X"84",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"d8",X"03",X"b2",X"03",X"19",X"03",X"b2",X"d8",X"03",X"b2",X"19",X"03",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"2e",X"ed",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"51",X"18",X"8e",X"8e",X"8e",X"8e",X"18",X"24",X"8e",X"8e",X"8e",X"8e",X"8e",X"18",X"41",X"a1",X"f5",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"06",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"0b",X"1b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"ed",X"03",X"75",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"b2",X"2e",X"00",X"1b",X"15",X"51",X"51",X"51",X"15",X"15",X"51",X"15",X"62",X"51",X"62",X"62",X"62",X"f5",X"f5",X"3d",X"cf",X"e9",X"62",X"1b",X"0b",X"00",X"0b",X"3c",X"0b",X"2e",X"03",X"1a",X"03",X"2e",X"0b",X"3c",X"0b",X"0b",X"25",X"4d",X"4d",X"4d",X"e9",X"4d",X"4d",X"4d",X"4d",X"3d",X"4d",X"ea",X"19",X"42",X"19",X"42",X"19",X"ea",X"bf",X"ea",X"75",X"19",X"75",X"75",X"0b",X"1b",X"19",X"75",X"75",X"19",X"0b",X"00",X"0b",X"1b",X"0b",X"2e",X"75",X"03",X"b2",X"03",X"03",X"03",X"b2",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"b2",X"27",X"03",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"f4",X"70",X"f3",X"82",X"70",X"82",X"82",X"70",X"82",X"82",X"70",X"82",X"82",X"4a",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"3f",X"6d",X"f0",X"7c",X"9e",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"b2",X"19",X"03",X"03",X"b2",X"19",X"71",X"19",X"71",X"03",X"b2",X"03",X"03",X"1a",X"03",X"2e",X"2f",X"62",X"62",X"15",X"cf",X"62",X"51",X"62",X"51",X"51",X"0f",X"51",X"f5",X"8e",X"8e",X"8e",X"8e",X"18",X"8e",X"a1",X"51",X"a1",X"51",X"51",X"15",X"f5",X"51",X"62",X"15",X"f5",X"51",X"62",X"ed",X"2e",X"03",X"75",X"03",X"b2",X"d8",X"75",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"0b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"7c",X"aa",X"aa",X"84",X"0b",X"1b",X"0b",X"79",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"d8",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"4d",X"0b",X"0b",X"3a",X"51",X"15",X"3a",X"51",X"51",X"62",X"62",X"cf",X"15",X"f5",X"62",X"cf",X"3d",X"cf",X"3d",X"3d",X"3d",X"3d",X"cf",X"e4",X"0b",X"0b",X"0b",X"3c",X"0b",X"2e",X"03",X"1a",X"03",X"2e",X"19",X"0b",X"1b",X"0b",X"3a",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"42",X"ea",X"19",X"ea",X"ea",X"75",X"ea",X"19",X"75",X"19",X"1a",X"19",X"3c",X"0b",X"75",X"75",X"19",X"75",X"b2",X"0b",X"0b",X"00",X"0b",X"2e",X"75",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"19",X"b2",X"19",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"82",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5d",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"9e",X"aa",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"27",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"75",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"2e",X"54",X"62",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"cf",X"15",X"62",X"a1",X"18",X"18",X"24",X"18",X"45",X"8e",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"15",X"f5",X"cf",X"15",X"62",X"51",X"f0",X"e5",X"03",X"b2",X"03",X"19",X"b2",X"27",X"03",X"1a",X"03",X"b2",X"27",X"03",X"b2",X"19",X"b2",X"19",X"71",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"3c",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"7c",X"9e",X"98",X"0b",X"0b",X"1b",X"2f",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"19",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"2e",X"1b",X"0b",X"3a",X"15",X"51",X"15",X"51",X"51",X"15",X"51",X"62",X"15",X"62",X"62",X"f5",X"3d",X"3d",X"cf",X"3d",X"3d",X"3d",X"5d",X"00",X"0b",X"3c",X"0b",X"3c",X"0b",X"2e",X"03",X"1a",X"03",X"2e",X"4d",X"3c",X"0b",X"00",X"0b",X"4d",X"4d",X"4d",X"4d",X"e9",X"4d",X"bf",X"4d",X"19",X"ea",X"ea",X"ea",X"42",X"19",X"42",X"75",X"ea",X"75",X"75",X"19",X"75",X"0b",X"00",X"75",X"19",X"75",X"19",X"b2",X"1b",X"0b",X"0b",X"3c",X"ec",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"19",X"b2",X"03",X"03",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"92",X"aa",X"84",X"0b",X"0b",X"1b",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"19",X"71",X"19",X"71",X"19",X"71",X"19",X"03",X"b2",X"27",X"19",X"03",X"cc",X"2f",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"51",X"18",X"24",X"18",X"18",X"18",X"8e",X"0f",X"62",X"15",X"cf",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"ed",X"2e",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"27",X"19",X"71",X"19",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"27",X"0b",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"1b",X"83",X"2f",X"03",X"b2",X"03",X"1a",X"71",X"19",X"71",X"19",X"71",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"03",X"03",X"b2",X"03",X"03",X"03",X"75",X"03",X"b2",X"4d",X"3c",X"0b",X"51",X"15",X"3a",X"51",X"15",X"62",X"62",X"62",X"62",X"cf",X"62",X"cf",X"3d",X"cf",X"3d",X"25",X"3d",X"3d",X"3d",X"62",X"1b",X"1b",X"0b",X"0b",X"0b",X"3c",X"0b",X"2e",X"03",X"b2",X"03",X"cc",X"2e",X"0b",X"0b",X"00",X"0b",X"4d",X"4d",X"4d",X"4d",X"4d",X"4d",X"3d",X"4d",X"ea",X"ea",X"ea",X"ea",X"ea",X"19",X"ea",X"19",X"75",X"19",X"75",X"19",X"1b",X"0b",X"19",X"75",X"75",X"19",X"1a",X"1b",X"0b",X"3c",X"3c",X"25",X"4d",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"3b",X"6d",X"f0",X"3f",X"6d",X"aa",X"9e",X"aa",X"aa",X"98",X"1b",X"0b",X"0b",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"19",X"71",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"2e",X"ed",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"15",X"f5",X"62",X"62",X"f5",X"18",X"18",X"24",X"18",X"24",X"18",X"0f",X"62",X"51",X"62",X"62",X"15",X"cf",X"15",X"51",X"62",X"15",X"51",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"71",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"75",X"03",X"03",X"19",X"71",X"19",X"03",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"b2",X"1b",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"60",X"ba",X"0b",X"0b",X"0b",X"2f",X"19",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"27",X"19",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"19",X"71",X"19",X"03",X"4d",X"2e",X"1b",X"3c",X"3a",X"51",X"15",X"51",X"15",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"f5",X"3d",X"cf",X"3d",X"3d",X"3d",X"3d",X"cf",X"17",X"1b",X"3c",X"0b",X"3c",X"0b",X"3c",X"2e",X"03",X"1a",X"03",X"03",X"cc",X"1b",X"0b",X"00",X"0b",X"4d",X"4d",X"4d",X"73",X"19",X"4d",X"fc",X"bf",X"ea",X"ea",X"19",X"ea",X"ea",X"75",X"ea",X"75",X"19",X"75",X"aa",X"75",X"e4",X"75",X"75",X"19",X"75",X"b2",X"0b",X"00",X"0b",X"0b",X"3d",X"e9",X"19",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"6d",X"aa",X"7c",X"aa",X"60",X"98",X"0b",X"0b",X"1b",X"03",X"1a",X"03",X"b2",X"19",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"19",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"2e",X"2f",X"62",X"62",X"15",X"cf",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"a1",X"18",X"8f",X"18",X"5b",X"18",X"8e",X"0f",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"62",X"cf",X"62",X"2f",X"2e",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"06",X"03",X"03",X"1a",X"03",X"19",X"71",X"19",X"71",X"03",X"1a",X"71",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"03",X"03",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",
    X"9e",X"aa",X"9e",X"aa",X"98",X"0b",X"1b",X"0b",X"79",X"03",X"b2",X"03",X"03",X"b2",X"19",X"71",X"19",X"03",X"b2",X"27",X"75",X"03",X"75",X"03",X"71",X"03",X"75",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"03",X"e5",X"03",X"1a",X"4d",X"3c",X"0b",X"51",X"15",X"51",X"15",X"51",X"62",X"62",X"15",X"62",X"62",X"cf",X"3d",X"cf",X"3d",X"3d",X"25",X"3d",X"3d",X"3d",X"3d",X"cf",X"0b",X"0b",X"3c",X"0b",X"0b",X"2e",X"03",X"1a",X"03",X"03",X"1a",X"03",X"2e",X"1b",X"0b",X"0b",X"3c",X"4d",X"4d",X"4d",X"4d",X"42",X"4d",X"fc",X"19",X"42",X"ea",X"ea",X"bf",X"ea",X"75",X"19",X"75",X"75",X"19",X"75",X"19",X"1a",X"19",X"75",X"75",X"1a",X"1b",X"0b",X"1b",X"0b",X"4d",X"3d",X"27",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"b2",X"19",X"03",X"03",X"b2",X"03",X"03",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"79",X"6d",X"f0",X"3f",X"aa",X"9e",X"aa",X"aa",X"23",X"0b",X"1b",X"0b",X"19",X"03",X"75",X"03",X"b2",X"03",X"1a",X"b2",X"27",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"71",X"19",X"b2",X"27",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"19",X"b2",X"27",X"75",X"2e",X"54",X"62",X"51",X"62",X"15",X"62",X"cf",X"62",X"51",X"62",X"51",X"62",X"f5",X"24",X"18",X"5b",X"18",X"8f",X"18",X"f5",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"61",X"2e",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"19",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"1b",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"ed",X"03",X"19",X"03",X"1a",X"03",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"1a",X"ec",X"1b",X"2e",X"03",X"4d",X"2e",X"3c",X"0b",X"3a",X"51",X"15",X"51",X"15",X"62",X"51",X"62",X"3a",X"f5",X"62",X"f5",X"3d",X"cf",X"3d",X"3d",X"3d",X"3d",X"3d",X"3d",X"62",X"3c",X"0b",X"0b",X"ec",X"03",X"1a",X"03",X"71",X"19",X"b2",X"03",X"b2",X"2e",X"0b",X"3c",X"0b",X"3c",X"4d",X"4d",X"ea",X"4d",X"bf",X"ea",X"ea",X"ea",X"ea",X"ea",X"ea",X"75",X"ea",X"75",X"75",X"19",X"75",X"75",X"19",X"75",X"19",X"75",X"19",X"b2",X"0b",X"00",X"0b",X"1b",X"4d",X"e9",X"19",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"00",X"00",X"fb",X"00",X"a4",X"91",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"4f",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"6d",X"aa",X"7c",X"aa",X"9e",X"98",X"0b",X"0b",X"0b",X"d8",X"b2",X"03",X"03",X"03",X"75",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"03",X"b2",X"03",X"cc",X"2f",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"15",X"62",X"62",X"51",X"f5",X"18",X"5b",X"18",X"30",X"18",X"8e",X"34",X"51",X"62",X"62",X"cf",X"15",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"71",X"19",X"b2",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"03",X"19",X"0b",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"28",X"03",X"b2",X"03",X"03",X"b2",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"19",X"71",X"19",X"03",X"2e",X"0b",X"2e",X"03",X"1a",X"2e",X"3c",X"0b",X"3c",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"00",X"0b",X"0b",X"1b",X"0b",X"0b",X"00",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"2e",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"ec",X"0b",X"1b",X"0b",X"00",X"ea",X"4d",X"ea",X"4d",X"42",X"bf",X"ea",X"ea",X"ea",X"19",X"ea",X"19",X"75",X"19",X"75",X"19",X"75",X"75",X"19",X"1a",X"75",X"19",X"1a",X"1b",X"0b",X"0b",X"00",X"75",X"2e",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"f4",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"9e",X"aa",X"2c",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"b2",X"19",X"71",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"03",X"2e",X"2f",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"cf",X"62",X"51",X"62",X"f5",X"24",X"18",X"30",X"24",X"c7",X"18",X"41",X"62",X"62",X"51",X"62",X"62",X"62",X"cf",X"62",X"51",X"62",X"51",X"62",X"ed",X"2e",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"75",X"03",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"71",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"0b",X"1b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"33",X"0b",X"0b",X"0b",X"79",X"1a",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"71",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"2e",X"3c",X"0b",X"2e",X"03",X"03",X"cc",X"3c",X"0b",X"1b",X"0b",X"3c",X"0b",X"1b",X"3c",X"1b",X"0b",X"3c",X"1b",X"3c",X"0b",X"1b",X"0b",X"00",X"0b",X"0b",X"1b",X"0b",X"3c",X"0b",X"2e",X"03",X"1a",X"03",X"b2",X"03",X"75",X"03",X"19",X"b2",X"27",X"19",X"1a",X"2e",X"3c",X"0b",X"0b",X"0b",X"19",X"4d",X"19",X"ea",X"ea",X"ea",X"bf",X"ea",X"ea",X"75",X"ea",X"75",X"19",X"75",X"75",X"19",X"1a",X"19",X"75",X"19",X"75",X"b2",X"1b",X"0b",X"3c",X"0b",X"19",X"2e",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"12",X"aa",X"92",X"61",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"b2",X"03",X"03",X"b2",X"27",X"19",X"71",X"19",X"71",X"19",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"21",X"54",X"62",X"62",X"15",X"cf",X"62",X"51",X"62",X"62",X"15",X"62",X"51",X"f5",X"18",X"8f",X"c7",X"18",X"30",X"18",X"a9",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"15",X"62",X"62",X"15",X"62",X"61",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"1a",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"7c",X"9e",X"98",X"0b",X"1b",X"0b",X"2f",X"03",X"03",X"b2",X"03",X"b2",X"d8",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"19",X"71",X"19",X"71",X"19",X"71",X"19",X"03",X"03",X"1a",X"03",X"03",X"19",X"ec",X"0b",X"1b",X"2e",X"03",X"1a",X"03",X"2e",X"2e",X"ec",X"2e",X"2e",X"ec",X"2e",X"2e",X"2e",X"2e",X"3c",X"0b",X"e9",X"30",X"cc",X"2e",X"2e",X"2e",X"ec",X"cc",X"cc",X"2e",X"ec",X"27",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"cc",X"19",X"1b",X"0b",X"00",X"0b",X"4d",X"ea",X"ea",X"ea",X"ea",X"ea",X"19",X"ea",X"75",X"19",X"1a",X"75",X"19",X"75",X"19",X"75",X"75",X"19",X"75",X"b2",X"0b",X"0b",X"3c",X"0b",X"75",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"19",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"00",X"00",X"f4",X"3c",X"a4",X"91",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"f4",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"2c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"d8",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"2e",X"ed",X"62",X"51",X"62",X"62",X"62",X"15",X"51",X"f5",X"51",X"62",X"15",X"41",X"8e",X"a4",X"8f",X"30",X"8f",X"18",X"41",X"62",X"15",X"62",X"51",X"62",X"15",X"62",X"62",X"cf",X"62",X"51",X"62",X"ed",X"2e",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"75",X"03",X"71",X"19",X"71",X"03",X"1a",X"03",X"19",X"03",X"b2",X"19",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"0b",X"0b",X"1b",X"17",X"f0",X"6d",X"3f",X"54",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"2f",X"03",X"1a",X"03",X"03",X"19",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"27",X"19",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"19",X"71",X"19",X"71",X"2e",X"0b",X"00",X"2e",X"0b",X"2e",X"03",X"1a",X"03",X"19",X"b2",X"19",X"71",X"19",X"03",X"1a",X"ec",X"0b",X"0b",X"3d",X"03",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"2e",X"4d",X"1b",X"0b",X"0b",X"3c",X"ea",X"ea",X"ea",X"ea",X"ea",X"bf",X"75",X"ea",X"19",X"75",X"19",X"75",X"75",X"19",X"1a",X"19",X"75",X"75",X"19",X"0b",X"3c",X"0b",X"0b",X"75",X"2e",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"00",X"00",X"fb",X"00",X"8f",X"fb",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"ad",X"0b",X"33",X"6d",X"3f",X"6d",X"3f",X"aa",X"9e",X"aa",X"9e",X"98",X"1b",X"0b",X"0b",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"03",X"1a",X"2e",X"2f",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"f5",X"62",X"62",X"f5",X"18",X"c7",X"c7",X"c7",X"c7",X"45",X"41",X"51",X"62",X"62",X"62",X"cf",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"19",X"03",X"b2",X"19",X"71",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"7c",X"aa",X"9e",X"98",X"1b",X"83",X"0b",X"2f",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"75",X"03",X"b2",X"03",X"03",X"19",X"71",X"75",X"71",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"2e",X"1b",X"0b",X"2e",X"00",X"1b",X"2e",X"03",X"b2",X"03",X"03",X"03",X"19",X"03",X"b2",X"03",X"2e",X"19",X"3c",X"4d",X"19",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"19",X"b2",X"03",X"2e",X"2e",X"2e",X"2e",X"3c",X"0b",X"00",X"0b",X"19",X"ea",X"ea",X"ea",X"19",X"ea",X"75",X"75",X"19",X"75",X"75",X"19",X"75",X"19",X"75",X"75",X"19",X"75",X"1b",X"0b",X"3c",X"0b",X"1b",X"2e",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"00",X"00",X"f4",X"3c",X"a4",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"3b",X"f0",X"6d",X"f0",X"6d",X"aa",X"7c",X"aa",X"7c",X"61",X"0b",X"0b",X"1b",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"75",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"2e",X"ed",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"cf",X"15",X"62",X"51",X"41",X"8e",X"8e",X"8e",X"8e",X"18",X"8e",X"41",X"62",X"62",X"51",X"15",X"51",X"62",X"51",X"62",X"51",X"62",X"cf",X"15",X"98",X"2e",X"03",X"19",X"03",X"b2",X"19",X"03",X"b2",X"03",X"b2",X"19",X"03",X"03",X"19",X"b2",X"27",X"19",X"03",X"b2",X"03",X"75",X"03",X"03",X"b2",X"27",X"75",X"03",X"b2",X"03",X"1a",X"03",X"71",X"19",X"03",X"19",X"0b",X"3c",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"9e",X"2c",X"ba",X"0b",X"1b",X"0b",X"79",X"03",X"71",X"19",X"03",X"19",X"03",X"b2",X"19",X"03",X"b2",X"03",X"27",X"19",X"71",X"19",X"71",X"19",X"03",X"03",X"19",X"71",X"19",X"03",X"b2",X"27",X"1a",X"03",X"03",X"21",X"0b",X"3c",X"2e",X"1b",X"0b",X"2e",X"03",X"19",X"21",X"2e",X"2e",X"ec",X"2e",X"03",X"19",X"21",X"75",X"0b",X"4d",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"2e",X"03",X"1a",X"03",X"19",X"03",X"19",X"03",X"03",X"03",X"f2",X"2e",X"3c",X"2e",X"83",X"2e",X"1b",X"0b",X"0b",X"0b",X"19",X"ea",X"ea",X"ea",X"19",X"ea",X"75",X"19",X"75",X"19",X"75",X"75",X"19",X"75",X"19",X"75",X"75",X"3c",X"0b",X"0b",X"3c",X"0b",X"ec",X"27",X"19",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"75",X"03",X"1a",X"03",X"00",X"00",X"fb",X"00",X"a4",X"91",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",X"9e",X"aa",X"9e",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"71",X"03",X"19",X"03",X"1a",X"03",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"03",X"21",X"f0",X"62",X"15",X"62",X"cf",X"62",X"62",X"15",X"f5",X"51",X"62",X"62",X"41",X"41",X"f5",X"41",X"41",X"34",X"f5",X"41",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"ed",X"2e",X"03",X"b2",X"27",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"71",X"19",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"75",X"03",X"b2",X"03",X"0b",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"2f",X"03",X"1a",X"03",X"b2",X"27",X"1a",X"03",X"03",X"b2",X"03",X"19",X"b2",X"27",X"19",X"03",X"1a",X"03",X"03",X"1a",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"2e",X"1b",X"0b",X"2e",X"0b",X"3c",X"2e",X"2e",X"2e",X"1b",X"0b",X"0b",X"0b",X"3c",X"2e",X"2e",X"03",X"4d",X"1b",X"75",X"2e",X"03",X"1a",X"03",X"b2",X"03",X"03",X"75",X"03",X"1a",X"03",X"1a",X"ec",X"0b",X"2e",X"2e",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"47",X"db",X"ec",X"0b",X"1b",X"2e",X"ad",X"2e",X"1b",X"0b",X"3c",X"0b",X"19",X"ea",X"75",X"ea",X"75",X"19",X"75",X"19",X"75",X"75",X"19",X"1a",X"75",X"19",X"1a",X"19",X"1b",X"0b",X"3c",X"0b",X"0b",X"2e",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"19",X"71",X"27",X"03",X"b2",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"7c",X"aa",X"9e",X"98",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"b2",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"2e",X"54",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"62",X"cf",X"15",X"f5",X"51",X"62",X"15",X"51",X"62",X"51",X"62",X"15",X"62",X"61",X"2e",X"03",X"75",X"03",X"b2",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"75",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"19",X"71",X"19",X"71",X"19",X"03",X"75",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"92",X"61",X"0b",X"0b",X"83",X"2f",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"27",X"19",X"03",X"03",X"1a",X"03",X"2e",X"3c",X"0b",X"2e",X"3c",X"0b",X"2e",X"1b",X"0b",X"3c",X"1b",X"0b",X"3c",X"0b",X"00",X"0b",X"2e",X"4d",X"00",X"75",X"2e",X"2e",X"03",X"1a",X"03",X"19",X"b2",X"03",X"03",X"03",X"e5",X"03",X"2e",X"00",X"2e",X"0b",X"2e",X"19",X"03",X"19",X"03",X"e8",X"9c",X"db",X"2e",X"0b",X"00",X"2e",X"e2",X"07",X"2e",X"3c",X"0b",X"0b",X"0b",X"19",X"ea",X"19",X"ea",X"75",X"75",X"19",X"75",X"19",X"1a",X"19",X"19",X"1a",X"19",X"75",X"0b",X"3c",X"0b",X"0b",X"3c",X"2e",X"03",X"19",X"03",X"71",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"75",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"9e",X"aa",X"2c",X"aa",X"33",X"0b",X"1b",X"0b",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"27",X"75",X"03",X"b2",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"19",X"2e",X"2f",X"62",X"62",X"62",X"62",X"15",X"62",X"62",X"15",X"cf",X"15",X"62",X"15",X"62",X"62",X"15",X"cf",X"15",X"62",X"51",X"62",X"62",X"62",X"15",X"cf",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"ed",X"2e",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"71",X"19",X"03",X"19",X"71",X"19",X"71",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"27",X"19",X"03",X"75",X"03",X"b2",X"03",X"0b",X"0b",X"1b",X"33",X"f0",X"6d",X"3f",X"6d",
    X"aa",X"7c",X"0d",X"aa",X"98",X"0b",X"1b",X"0b",X"2f",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"d8",X"75",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"b2",X"03",X"1a",X"ec",X"0b",X"1b",X"2e",X"1b",X"0b",X"0b",X"3c",X"0b",X"1b",X"0b",X"0b",X"3c",X"0b",X"0b",X"00",X"1b",X"e9",X"1b",X"19",X"2e",X"06",X"2e",X"03",X"03",X"b2",X"03",X"19",X"b2",X"2e",X"1b",X"2e",X"2e",X"1b",X"0b",X"00",X"2e",X"03",X"b2",X"27",X"b5",X"3e",X"10",X"e2",X"2e",X"1b",X"0b",X"2e",X"b5",X"3e",X"b5",X"2e",X"1b",X"0b",X"3c",X"0b",X"75",X"ea",X"75",X"75",X"19",X"75",X"75",X"75",X"19",X"75",X"75",X"75",X"19",X"75",X"3c",X"1b",X"0b",X"3c",X"0b",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"82",X"3c",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"70",X"f4",X"4f",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"9e",X"aa",X"7c",X"61",X"0b",X"0b",X"1b",X"03",X"1a",X"03",X"b2",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"cc",X"2f",X"62",X"51",X"62",X"15",X"cf",X"62",X"51",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"cf",X"62",X"62",X"51",X"62",X"ed",X"2e",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"19",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"1a",X"e4",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"7c",X"aa",X"61",X"0b",X"1b",X"0b",X"79",X"03",X"19",X"03",X"b2",X"27",X"75",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"2e",X"0b",X"3c",X"2e",X"3c",X"0b",X"3c",X"0b",X"8b",X"f3",X"f3",X"ae",X"8b",X"0b",X"1b",X"0b",X"0b",X"3d",X"1b",X"1a",X"2e",X"19",X"0b",X"2e",X"1a",X"03",X"03",X"b2",X"03",X"2e",X"3c",X"2e",X"2e",X"0b",X"3c",X"0b",X"30",X"03",X"1a",X"e2",X"3e",X"3e",X"b5",X"9c",X"2e",X"3c",X"0b",X"2e",X"47",X"3e",X"b5",X"e2",X"2e",X"3c",X"0b",X"0b",X"1b",X"0b",X"75",X"19",X"75",X"75",X"19",X"75",X"19",X"75",X"19",X"75",X"19",X"1a",X"1b",X"0b",X"0b",X"0b",X"3c",X"2e",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"00",X"00",X"fb",X"00",X"a4",X"4f",X"82",X"70",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"82",X"82",X"f4",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"3b",X"6d",X"f0",X"6d",X"f0",X"7c",X"aa",X"9e",X"aa",X"74",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"19",X"03",X"b2",X"19",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"03",X"2e",X"54",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"15",X"62",X"51",X"62",X"15",X"62",X"62",X"62",X"15",X"62",X"51",X"15",X"62",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"27",X"75",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"19",X"3c",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"9e",X"aa",X"60",X"98",X"0b",X"0b",X"0b",X"2f",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"19",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"2e",X"3c",X"0b",X"2e",X"1b",X"1b",X"0b",X"4e",X"f3",X"f3",X"ae",X"82",X"ae",X"ae",X"8b",X"0b",X"3c",X"2e",X"0b",X"1a",X"ec",X"bf",X"00",X"2e",X"03",X"03",X"1a",X"03",X"03",X"cc",X"1b",X"2e",X"2e",X"3c",X"0b",X"0b",X"2e",X"03",X"03",X"b5",X"3e",X"b5",X"3e",X"db",X"2e",X"1b",X"3c",X"2e",X"e2",X"10",X"47",X"83",X"0b",X"2e",X"1b",X"00",X"0b",X"3c",X"0b",X"75",X"19",X"75",X"75",X"19",X"75",X"75",X"75",X"19",X"75",X"19",X"0b",X"3c",X"0b",X"3c",X"0b",X"2e",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"00",X"00",X"f4",X"3c",X"8f",X"4f",X"f4",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"4a",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"9e",X"aa",X"7c",X"aa",X"98",X"0b",X"0b",X"0b",X"75",X"03",X"71",X"19",X"71",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"19",X"b2",X"27",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"27",X"1a",X"03",X"03",X"1a",X"03",X"03",X"71",X"03",X"1a",X"03",X"2e",X"ed",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"62",X"62",X"cf",X"15",X"f5",X"51",X"62",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"cf",X"62",X"2f",X"2e",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"03",X"75",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"71",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"0b",X"1b",X"0b",X"17",X"6d",X"3f",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"aa",X"ba",X"0b",X"0b",X"1b",X"61",X"03",X"75",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"27",X"19",X"03",X"b2",X"27",X"1a",X"03",X"03",X"19",X"03",X"2e",X"0b",X"0b",X"2e",X"b2",X"0b",X"0b",X"f3",X"8b",X"22",X"f3",X"ae",X"70",X"ae",X"39",X"ae",X"1b",X"2e",X"1b",X"1b",X"2e",X"4d",X"1b",X"30",X"03",X"1a",X"03",X"b2",X"19",X"2e",X"00",X"2e",X"2e",X"1b",X"0b",X"1b",X"2e",X"1b",X"66",X"07",X"3e",X"e2",X"10",X"e2",X"2e",X"1a",X"1b",X"2e",X"47",X"10",X"b5",X"83",X"0b",X"00",X"2e",X"19",X"1b",X"0b",X"1b",X"0b",X"75",X"19",X"75",X"75",X"19",X"75",X"19",X"75",X"75",X"75",X"1b",X"0b",X"00",X"0b",X"00",X"2e",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"00",X"00",X"fb",X"00",X"a4",X"4f",X"f4",X"fb",X"f4",X"4f",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"91",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"9e",X"aa",X"9e",X"98",X"0b",X"0b",X"1b",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"27",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"ec",X"f0",X"62",X"15",X"62",X"cf",X"62",X"15",X"62",X"cf",X"62",X"62",X"51",X"62",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"cf",X"62",X"15",X"f5",X"62",X"62",X"62",X"62",X"51",X"15",X"f5",X"ed",X"2e",X"19",X"b2",X"27",X"19",X"71",X"19",X"03",X"03",X"19",X"03",X"19",X"71",X"19",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"0b",X"0b",X"3c",X"33",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"9e",X"2c",X"61",X"0b",X"1b",X"0b",X"2f",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"1a",X"b2",X"27",X"30",X"3c",X"0b",X"ec",X"1a",X"3c",X"65",X"4e",X"f3",X"f3",X"ae",X"f3",X"ae",X"82",X"ae",X"39",X"8b",X"2e",X"b2",X"1b",X"3d",X"4d",X"1b",X"25",X"ec",X"03",X"19",X"03",X"03",X"e5",X"1b",X"2e",X"2e",X"00",X"0b",X"00",X"3d",X"cd",X"9c",X"3e",X"b5",X"db",X"e2",X"0b",X"2e",X"b2",X"0b",X"2e",X"e2",X"10",X"47",X"56",X"0b",X"2e",X"0b",X"2e",X"4d",X"1b",X"3c",X"0b",X"0b",X"75",X"19",X"75",X"75",X"19",X"75",X"19",X"75",X"19",X"3c",X"0b",X"0b",X"0b",X"0b",X"2e",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"00",X"00",X"f4",X"3c",X"8f",X"4f",X"f4",X"91",X"f4",X"f4",X"fb",X"fb",X"f4",X"fb",X"f4",X"4f",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",X"7c",X"aa",X"7c",X"aa",X"84",X"0b",X"1b",X"0b",X"d8",X"1a",X"03",X"b2",X"19",X"71",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"2e",X"98",X"51",X"62",X"62",X"15",X"51",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"cf",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"cf",X"62",X"15",X"cf",X"62",X"51",X"62",X"62",X"62",X"ed",X"2e",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"b2",X"27",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"0b",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"aa",X"ba",X"0b",X"0b",X"0b",X"77",X"03",X"19",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"2e",X"1b",X"0b",X"2e",X"1a",X"1b",X"8b",X"f3",X"6f",X"f3",X"f3",X"ae",X"82",X"ae",X"39",X"ae",X"39",X"2e",X"1a",X"3c",X"25",X"e9",X"3c",X"4d",X"2e",X"2e",X"2e",X"2e",X"ec",X"2e",X"0b",X"2e",X"ec",X"0b",X"1b",X"0b",X"25",X"1b",X"db",X"db",X"47",X"10",X"0b",X"e2",X"2e",X"1a",X"3c",X"2e",X"83",X"83",X"47",X"a3",X"0b",X"2e",X"ec",X"a3",X"25",X"ec",X"0b",X"1b",X"0b",X"00",X"75",X"19",X"75",X"75",X"75",X"19",X"75",X"75",X"0b",X"1b",X"0b",X"3c",X"1b",X"2e",X"03",X"b2",X"03",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"1a",X"00",X"00",X"fb",X"00",X"a4",X"4f",X"f4",X"fb",X"f4",X"91",X"f4",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"fb",X"f4",X"fb",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"9e",X"aa",X"9e",X"aa",X"98",X"0b",X"0b",X"0b",X"19",X"71",X"19",X"03",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"2e",X"2f",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"62",X"15",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"ed",X"2e",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"9e",X"aa",X"60",X"98",X"0b",X"1b",X"0b",X"28",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"19",X"71",X"19",X"71",X"03",X"1a",X"03",X"19",X"71",X"19",X"b2",X"2e",X"54",X"3c",X"2e",X"aa",X"0b",X"4e",X"8b",X"f3",X"22",X"ae",X"f3",X"ae",X"ae",X"ae",X"39",X"4a",X"39",X"6f",X"1b",X"32",X"d6",X"0b",X"3f",X"2e",X"2e",X"1b",X"0b",X"0b",X"2e",X"3c",X"2e",X"2e",X"0b",X"3c",X"0b",X"ea",X"d6",X"e2",X"b5",X"47",X"b5",X"1b",X"66",X"2e",X"aa",X"0b",X"2e",X"e2",X"0b",X"56",X"83",X"0b",X"2e",X"0b",X"2e",X"1b",X"e2",X"2e",X"0b",X"3c",X"0b",X"0b",X"75",X"19",X"75",X"19",X"75",X"19",X"75",X"3c",X"0b",X"3c",X"0b",X"0b",X"2e",X"03",X"19",X"03",X"19",X"b2",X"27",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"fb",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"7c",X"aa",X"61",X"0b",X"1b",X"0b",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"b2",X"27",X"19",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"19",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"03",X"2e",X"ed",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"cf",X"62",X"15",X"62",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"cf",X"62",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"cf",X"15",X"62",X"15",X"61",X"2e",X"03",X"19",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"75",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"19",X"b2",X"19",X"71",X"19",X"03",X"1a",X"1b",X"0b",X"0b",X"53",X"6d",X"f0",X"3f",X"6d",
    X"aa",X"7c",X"0d",X"aa",X"98",X"0b",X"1b",X"0b",X"79",X"1a",X"03",X"19",X"03",X"71",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"2e",X"2f",X"0b",X"2e",X"aa",X"0b",X"eb",X"f3",X"4e",X"f3",X"f3",X"ae",X"82",X"ae",X"39",X"ae",X"39",X"d1",X"65",X"0b",X"e9",X"32",X"0b",X"f0",X"6d",X"00",X"0b",X"3c",X"1b",X"2e",X"1b",X"2e",X"2e",X"00",X"0b",X"00",X"42",X"d6",X"2e",X"2e",X"83",X"0b",X"3c",X"83",X"2e",X"aa",X"0b",X"2e",X"b5",X"ad",X"0b",X"ad",X"1b",X"2e",X"1b",X"0b",X"ec",X"66",X"47",X"2e",X"1b",X"0b",X"3c",X"0b",X"75",X"19",X"75",X"75",X"75",X"19",X"0b",X"00",X"0b",X"0b",X"3c",X"2e",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"1a",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"3c",X"00",X"f4",X"fb",X"fb",X"00",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"00",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"3f",X"6d",X"f0",X"7c",X"9e",X"aa",X"12",X"98",X"0b",X"0b",X"0b",X"19",X"71",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"27",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"b2",X"2e",X"2f",X"62",X"62",X"15",X"cf",X"62",X"15",X"62",X"15",X"62",X"cf",X"62",X"62",X"62",X"51",X"51",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"03",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"0b",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"7c",X"aa",X"61",X"0b",X"0b",X"0b",X"79",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"27",X"75",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"cc",X"54",X"0b",X"2e",X"fc",X"0b",X"af",X"8b",X"f3",X"f3",X"ae",X"f3",X"0b",X"00",X"82",X"39",X"39",X"4a",X"8b",X"3c",X"73",X"32",X"0b",X"1b",X"0b",X"0b",X"00",X"0b",X"0b",X"2e",X"3c",X"2e",X"2e",X"1b",X"0b",X"0b",X"aa",X"2e",X"2e",X"f0",X"2e",X"0b",X"1b",X"00",X"2e",X"9e",X"1b",X"2e",X"1b",X"83",X"b5",X"e2",X"66",X"2e",X"3c",X"0b",X"2e",X"83",X"b5",X"83",X"2e",X"3c",X"0b",X"0b",X"0b",X"75",X"19",X"75",X"19",X"75",X"1b",X"0b",X"0b",X"3c",X"0b",X"2e",X"19",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"06",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"00",X"00",X"f4",X"3c",X"8f",X"3c",X"82",X"70",X"3c",X"f4",X"00",X"2e",X"2e",X"2e",X"00",X"00",X"00",X"00",X"2e",X"2e",X"00",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"aa",X"2c",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"03",X"1a",X"03",X"1a",X"03",X"75",X"03",X"03",X"03",X"1a",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"2e",X"54",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"cf",X"62",X"62",X"62",X"62",X"51",X"62",X"15",X"f5",X"cf",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"f0",X"2e",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"b2",X"03",X"1a",X"03",X"0b",X"3c",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"9e",X"aa",X"60",X"98",X"0b",X"0b",X"1b",X"79",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"2e",X"aa",X"0b",X"d6",X"fc",X"0b",X"8b",X"46",X"eb",X"f3",X"f3",X"1b",X"0b",X"03",X"0b",X"82",X"d1",X"39",X"f3",X"0b",X"42",X"2e",X"3c",X"3c",X"0b",X"1b",X"0b",X"0b",X"1b",X"2e",X"0b",X"f3",X"2e",X"1b",X"0b",X"1b",X"9e",X"2e",X"ec",X"54",X"3c",X"2e",X"00",X"0b",X"2e",X"aa",X"0b",X"2e",X"56",X"83",X"0b",X"0b",X"1b",X"2e",X"1b",X"0b",X"2e",X"1b",X"56",X"0b",X"00",X"2e",X"1b",X"0b",X"00",X"0b",X"75",X"19",X"75",X"75",X"3c",X"0b",X"3c",X"0b",X"3c",X"2e",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"00",X"00",X"fb",X"00",X"a4",X"00",X"82",X"82",X"3c",X"00",X"00",X"2e",X"2e",X"00",X"f4",X"fb",X"fb",X"f4",X"3c",X"2e",X"00",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"12",X"aa",X"9e",X"54",X"1b",X"0b",X"0b",X"19",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"2e",X"2f",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"cf",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"cf",X"62",X"62",X"15",X"f5",X"cf",X"15",X"98",X"2e",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"84",X"0b",X"1b",X"0b",X"ed",X"03",X"19",X"03",X"75",X"03",X"b2",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"03",X"19",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"2e",X"aa",X"0b",X"d6",X"42",X"3c",X"eb",X"8b",X"f3",X"22",X"ae",X"0b",X"0b",X"03",X"1a",X"1b",X"39",X"39",X"ae",X"0b",X"f0",X"2e",X"0b",X"0b",X"0b",X"3c",X"0b",X"4a",X"39",X"2e",X"1b",X"ae",X"f3",X"6f",X"00",X"0b",X"2f",X"2e",X"2e",X"98",X"1b",X"2e",X"83",X"e2",X"2e",X"aa",X"0b",X"d6",X"83",X"0b",X"0b",X"0b",X"83",X"2e",X"0b",X"3c",X"2e",X"0b",X"1b",X"00",X"3c",X"3c",X"2e",X"7d",X"0b",X"3c",X"0b",X"0b",X"75",X"19",X"0b",X"00",X"0b",X"0b",X"0b",X"ec",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"00",X"00",X"f4",X"3c",X"8f",X"4f",X"3c",X"00",X"fb",X"00",X"2e",X"2e",X"2e",X"00",X"fb",X"f4",X"fb",X"f4",X"3c",X"2e",X"00",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7f",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"6d",X"aa",X"7c",X"aa",X"74",X"0b",X"0b",X"0b",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"03",X"19",X"03",X"1a",X"03",X"b2",X"d8",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"21",X"2f",X"f5",X"51",X"62",X"62",X"62",X"cf",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"15",X"51",X"62",X"62",X"51",X"62",X"62",X"ed",X"2e",X"03",X"75",X"03",X"b2",X"03",X"19",X"b2",X"03",X"b2",X"03",X"75",X"03",X"1a",X"03",X"03",X"b2",X"27",X"1a",X"03",X"75",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"0b",X"0b",X"1b",X"17",X"3f",X"6d",X"6d",X"f0",
    X"9e",X"aa",X"9e",X"7c",X"61",X"0b",X"0b",X"0b",X"28",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"71",X"19",X"19",X"b2",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"21",X"aa",X"1b",X"d6",X"4d",X"1b",X"8b",X"f3",X"4e",X"f3",X"f3",X"0b",X"1b",X"0b",X"0b",X"00",X"f3",X"4a",X"d1",X"0b",X"3c",X"2e",X"0b",X"1b",X"0b",X"d1",X"39",X"39",X"ae",X"2e",X"ad",X"f3",X"ae",X"8b",X"1b",X"0b",X"54",X"2e",X"2e",X"aa",X"0b",X"d6",X"2e",X"e2",X"2e",X"fc",X"0b",X"d6",X"50",X"0b",X"1b",X"83",X"66",X"2e",X"00",X"0b",X"2e",X"00",X"0b",X"0b",X"0b",X"e2",X"66",X"2e",X"7d",X"0b",X"0b",X"3c",X"0b",X"75",X"1b",X"0b",X"00",X"0b",X"1b",X"2e",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"71",X"19",X"71",X"19",X"03",X"00",X"00",X"fb",X"00",X"a4",X"4f",X"f4",X"fb",X"f4",X"3c",X"2e",X"2e",X"2e",X"00",X"00",X"00",X"00",X"00",X"00",X"2e",X"00",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"cd",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"9e",X"aa",X"98",X"1b",X"0b",X"0b",X"d8",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"19",X"b2",X"27",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"03",X"2e",X"54",X"15",X"62",X"62",X"51",X"62",X"15",X"62",X"15",X"f5",X"51",X"cf",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"15",X"62",X"61",X"2e",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"19",X"0b",X"3c",X"0b",X"33",X"6d",X"f0",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"79",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"71",X"27",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"03",X"b2",X"03",X"2e",X"ea",X"0b",X"4d",X"e9",X"00",X"af",X"6f",X"f3",X"f3",X"ae",X"f3",X"0b",X"1b",X"0b",X"1b",X"8b",X"39",X"d1",X"0b",X"1b",X"2e",X"3c",X"d1",X"ff",X"39",X"fb",X"39",X"d1",X"82",X"ae",X"82",X"f3",X"f3",X"3c",X"0b",X"ed",X"2e",X"2e",X"aa",X"0b",X"d6",X"2e",X"2e",X"ec",X"fc",X"0b",X"d6",X"b5",X"0b",X"56",X"b5",X"83",X"2e",X"1b",X"00",X"2e",X"0b",X"00",X"1b",X"0b",X"83",X"66",X"47",X"2e",X"2e",X"3c",X"0b",X"0b",X"00",X"0b",X"0b",X"3c",X"0b",X"3c",X"2e",X"03",X"b2",X"19",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"03",X"03",X"19",X"03",X"b2",X"03",X"00",X"00",X"f4",X"3c",X"8f",X"4f",X"f4",X"fb",X"f4",X"3c",X"2e",X"2e",X"2e",X"00",X"fb",X"f4",X"fb",X"f4",X"3c",X"2e",X"00",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"7c",X"9e",X"aa",X"33",X"0b",X"0b",X"1b",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"19",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"19",X"2e",X"ed",X"62",X"51",X"15",X"62",X"51",X"62",X"62",X"cf",X"15",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"cf",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"cf",X"15",X"62",X"62",X"51",X"2f",X"2e",X"03",X"19",X"03",X"b2",X"27",X"19",X"71",X"19",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"75",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"60",X"61",X"0b",X"0b",X"0b",X"2f",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"2e",X"fc",X"1b",X"73",X"4d",X"1b",X"0b",X"f3",X"4e",X"f3",X"f3",X"ae",X"ae",X"f3",X"48",X"4e",X"0b",X"4e",X"d1",X"0b",X"0b",X"2e",X"57",X"d1",X"39",X"d1",X"39",X"39",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"0b",X"0b",X"3c",X"2e",X"2e",X"aa",X"0b",X"e9",X"ec",X"0b",X"2e",X"4d",X"7f",X"d6",X"e2",X"83",X"83",X"3e",X"83",X"2e",X"1b",X"0b",X"2e",X"1b",X"00",X"0b",X"0b",X"56",X"83",X"83",X"0b",X"56",X"2e",X"1b",X"0b",X"0b",X"0b",X"00",X"0b",X"0b",X"2e",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"19",X"03",X"b2",X"19",X"71",X"19",X"b2",X"27",X"19",X"03",X"00",X"00",X"fb",X"00",X"a4",X"4f",X"f4",X"91",X"f4",X"3c",X"2e",X"2e",X"2e",X"00",X"f4",X"fb",X"f4",X"fb",X"00",X"2e",X"00",X"f4",X"3c",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"ad",X"1b",X"33",X"f0",X"6d",X"f0",X"6d",X"9e",X"aa",X"aa",X"7c",X"61",X"0b",X"1b",X"0b",X"03",X"b2",X"27",X"19",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"75",X"03",X"1a",X"03",X"75",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"03",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"03",X"2e",X"2f",X"62",X"62",X"62",X"cf",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"cf",X"62",X"62",X"51",X"15",X"f5",X"cf",X"62",X"15",X"cf",X"15",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"61",X"2e",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"06",X"03",X"b2",X"19",X"03",X"1a",X"03",X"71",X"19",X"1b",X"0b",X"0b",X"3b",X"6d",X"f0",X"3f",X"6d",
    X"aa",X"7c",X"0d",X"aa",X"98",X"0b",X"1b",X"0b",X"79",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"27",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"71",X"27",X"ec",X"fc",X"0b",X"4d",X"e9",X"3c",X"1b",X"8b",X"f3",X"f3",X"ae",X"f3",X"ae",X"82",X"ae",X"39",X"39",X"39",X"39",X"d1",X"1b",X"2e",X"d1",X"d1",X"d1",X"d1",X"39",X"4a",X"39",X"ae",X"ae",X"ae",X"f3",X"f3",X"0b",X"3c",X"0b",X"ec",X"2e",X"ea",X"3c",X"4d",X"2e",X"1b",X"2e",X"73",X"3c",X"4d",X"86",X"1b",X"96",X"10",X"83",X"2e",X"1a",X"3c",X"2e",X"0b",X"3c",X"1b",X"0b",X"56",X"83",X"e2",X"0b",X"83",X"03",X"21",X"2e",X"3c",X"1b",X"0b",X"2e",X"ec",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"03",X"19",X"03",X"71",X"19",X"b2",X"00",X"00",X"f4",X"3c",X"8f",X"4f",X"f4",X"fb",X"f4",X"00",X"2e",X"2e",X"2e",X"00",X"fb",X"f4",X"fb",X"f4",X"00",X"2e",X"00",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"7c",X"aa",X"9e",X"98",X"0b",X"0b",X"0b",X"03",X"1a",X"03",X"71",X"19",X"b2",X"27",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"19",X"b2",X"27",X"75",X"03",X"b2",X"27",X"19",X"03",X"b2",X"2e",X"f0",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"15",X"f5",X"51",X"62",X"62",X"62",X"15",X"51",X"f5",X"62",X"62",X"cf",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"2f",X"2e",X"1a",X"03",X"19",X"71",X"19",X"03",X"71",X"19",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"03",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"3c",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"7c",X"aa",X"61",X"0b",X"0b",X"0b",X"2f",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"d6",X"4d",X"1b",X"42",X"d6",X"0b",X"0b",X"f3",X"6f",X"f3",X"f3",X"ae",X"ae",X"82",X"d1",X"82",X"39",X"fb",X"d1",X"39",X"d1",X"d1",X"57",X"d1",X"39",X"d1",X"39",X"d1",X"82",X"39",X"ae",X"f3",X"ae",X"f3",X"1b",X"0b",X"0b",X"2e",X"2e",X"fc",X"0b",X"42",X"2e",X"3c",X"2e",X"d6",X"0b",X"e9",X"e9",X"1b",X"56",X"47",X"83",X"2e",X"b2",X"1b",X"2e",X"1b",X"00",X"0b",X"0b",X"e2",X"47",X"b5",X"0b",X"e8",X"03",X"1a",X"03",X"2e",X"0b",X"2e",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"75",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"00",X"00",X"fb",X"00",X"a4",X"4f",X"f4",X"fb",X"f4",X"00",X"2e",X"2e",X"2e",X"00",X"00",X"00",X"00",X"00",X"00",X"2e",X"00",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"9e",X"aa",X"2c",X"aa",X"98",X"0b",X"1b",X"0b",X"19",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"75",X"03",X"19",X"b2",X"19",X"03",X"1a",X"03",X"19",X"71",X"27",X"03",X"03",X"b2",X"03",X"03",X"19",X"b2",X"03",X"1a",X"03",X"21",X"f0",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"15",X"62",X"51",X"15",X"cf",X"62",X"15",X"79",X"2e",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"71",X"27",X"19",X"b2",X"27",X"19",X"03",X"b2",X"19",X"03",X"19",X"03",X"1a",X"03",X"b2",X"27",X"03",X"75",X"03",X"03",X"b2",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"79",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"d6",X"14",X"3c",X"fc",X"d6",X"0b",X"00",X"4e",X"f3",X"f3",X"ae",X"f3",X"ae",X"ae",X"82",X"39",X"d1",X"39",X"4a",X"57",X"d1",X"57",X"d1",X"d1",X"ff",X"39",X"4a",X"39",X"4a",X"ae",X"82",X"8b",X"3c",X"0b",X"0b",X"00",X"1b",X"2e",X"2e",X"ea",X"1b",X"ea",X"2e",X"1b",X"d6",X"d6",X"1b",X"ea",X"3d",X"5d",X"0b",X"56",X"47",X"2e",X"1a",X"1b",X"2e",X"00",X"0b",X"0b",X"1b",X"b5",X"47",X"0b",X"b5",X"e9",X"19",X"03",X"b2",X"27",X"30",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"03",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"75",X"03",X"19",X"03",X"1a",X"03",X"00",X"00",X"f4",X"3c",X"8f",X"4f",X"f4",X"fb",X"91",X"00",X"2e",X"2e",X"2e",X"00",X"fb",X"f4",X"fb",X"fb",X"00",X"2e",X"00",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"aa",X"12",X"aa",X"98",X"0b",X"0b",X"3c",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"71",X"03",X"03",X"1a",X"03",X"2e",X"1a",X"15",X"62",X"62",X"62",X"15",X"cf",X"15",X"51",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"cf",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"75",X"ec",X"03",X"1a",X"03",X"19",X"03",X"71",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"b2",X"27",X"19",X"03",X"b2",X"19",X"71",X"03",X"1a",X"03",X"0b",X"1b",X"0b",X"53",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"7c",X"aa",X"aa",X"84",X"0b",X"0b",X"1b",X"2f",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"fc",X"d6",X"0b",X"42",X"d6",X"1b",X"0b",X"0b",X"65",X"f3",X"f3",X"ae",X"82",X"70",X"d1",X"82",X"39",X"39",X"d1",X"d1",X"d1",X"d1",X"57",X"d1",X"39",X"d1",X"d1",X"39",X"ae",X"8b",X"0b",X"00",X"0b",X"0b",X"1b",X"0b",X"2e",X"db",X"ec",X"fc",X"0b",X"fc",X"2e",X"2f",X"73",X"ec",X"0b",X"42",X"e9",X"1b",X"0b",X"0b",X"56",X"2e",X"06",X"0b",X"2e",X"0b",X"0b",X"00",X"00",X"00",X"00",X"1a",X"03",X"3d",X"2e",X"03",X"75",X"03",X"71",X"75",X"03",X"19",X"03",X"b2",X"27",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"71",X"03",X"b2",X"03",X"03",X"b2",X"00",X"00",X"fb",X"00",X"a4",X"4f",X"f4",X"fb",X"f4",X"fb",X"00",X"2e",X"2e",X"00",X"fb",X"f4",X"fb",X"f4",X"3c",X"2e",X"00",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"60",X"aa",X"9e",X"aa",X"74",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"cc",X"1a",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"51",X"cf",X"15",X"62",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"cf",X"15",X"62",X"51",X"62",X"62",X"1a",X"2e",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"75",X"03",X"03",X"b2",X"03",X"19",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"19",X"0b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"9e",X"7c",X"61",X"0b",X"0b",X"83",X"2f",X"03",X"b2",X"27",X"19",X"03",X"b2",X"d8",X"03",X"1a",X"03",X"b2",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"ea",X"d6",X"0b",X"aa",X"2e",X"0b",X"3c",X"0b",X"1b",X"0b",X"ae",X"f3",X"ae",X"ae",X"ae",X"39",X"d1",X"4a",X"39",X"d1",X"ff",X"d1",X"57",X"d1",X"57",X"39",X"4a",X"39",X"0b",X"1b",X"0b",X"1b",X"0b",X"00",X"2e",X"2e",X"00",X"00",X"2e",X"e9",X"3c",X"42",X"2e",X"54",X"73",X"2e",X"3c",X"aa",X"2e",X"83",X"2e",X"1b",X"0b",X"2e",X"19",X"00",X"2e",X"1b",X"56",X"0b",X"00",X"00",X"00",X"03",X"03",X"2e",X"b2",X"30",X"03",X"2e",X"19",X"03",X"03",X"b2",X"d8",X"19",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"00",X"00",X"f4",X"3c",X"8f",X"4f",X"f4",X"fb",X"f4",X"fb",X"00",X"2e",X"2e",X"2e",X"00",X"00",X"00",X"00",X"2e",X"2e",X"00",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"7c",X"aa",X"98",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"b2",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"19",X"03",X"b2",X"19",X"71",X"27",X"1a",X"03",X"71",X"19",X"21",X"03",X"28",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"15",X"62",X"15",X"62",X"15",X"62",X"62",X"62",X"51",X"62",X"62",X"28",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"71",X"19",X"71",X"03",X"1a",X"03",X"b2",X"27",X"75",X"03",X"b2",X"03",X"0b",X"3c",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"2f",X"19",X"03",X"1a",X"71",X"19",X"03",X"1a",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"19",X"2e",X"00",X"aa",X"2e",X"0b",X"1b",X"0b",X"3c",X"0b",X"00",X"1b",X"65",X"ae",X"39",X"ae",X"39",X"39",X"d1",X"39",X"d1",X"d1",X"d1",X"d1",X"d1",X"d1",X"39",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"2e",X"ec",X"1b",X"00",X"0b",X"2e",X"4d",X"1b",X"1b",X"2e",X"aa",X"aa",X"2e",X"0b",X"54",X"2e",X"2e",X"b2",X"2e",X"e2",X"2e",X"75",X"1b",X"e9",X"56",X"e2",X"e2",X"0b",X"00",X"00",X"03",X"75",X"ec",X"1a",X"e9",X"ec",X"2e",X"2e",X"03",X"1a",X"03",X"b2",X"27",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"75",X"03",X"b2",X"03",X"00",X"00",X"fb",X"00",X"a4",X"4f",X"f4",X"fb",X"f4",X"91",X"f4",X"00",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"00",X"fb",X"f4",X"3c",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"cd",X"6d",X"f0",X"6d",X"3f",X"aa",X"60",X"aa",X"60",X"61",X"0b",X"0b",X"1b",X"d8",X"b2",X"03",X"19",X"b2",X"19",X"03",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"e5",X"03",X"1a",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"15",X"75",X"03",X"cc",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"0b",X"0b",X"0b",X"3b",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"9e",X"aa",X"60",X"61",X"0b",X"0b",X"0b",X"79",X"03",X"b2",X"03",X"03",X"19",X"b2",X"03",X"03",X"03",X"19",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"e5",X"0b",X"2f",X"2e",X"3c",X"0b",X"f3",X"0b",X"1b",X"0b",X"0b",X"0b",X"65",X"82",X"39",X"fb",X"39",X"d1",X"d1",X"57",X"d1",X"57",X"d1",X"d1",X"39",X"d1",X"39",X"ae",X"8b",X"0b",X"0b",X"1b",X"0b",X"2e",X"2e",X"2e",X"83",X"2e",X"d6",X"3c",X"0b",X"2e",X"aa",X"12",X"2e",X"3c",X"f0",X"2e",X"ec",X"1a",X"e4",X"2e",X"2e",X"19",X"0b",X"3d",X"50",X"b5",X"83",X"0b",X"00",X"03",X"b2",X"27",X"2e",X"1a",X"4d",X"2e",X"2e",X"06",X"2e",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"f4",X"fb",X"f4",X"3c",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"6d",X"36",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"75",X"03",X"19",X"b2",X"03",X"03",X"03",X"b2",X"2e",X"ec",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"2e",X"2e",X"03",X"b2",X"03",X"2e",X"03",X"1a",X"75",X"15",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"62",X"75",X"19",X"b2",X"2e",X"03",X"03",X"b2",X"2e",X"ec",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"2e",X"2e",X"ec",X"2e",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"0b",X"1b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"0d",X"aa",X"98",X"0b",X"1b",X"0b",X"2f",X"03",X"19",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"21",X"1b",X"54",X"2e",X"1b",X"0b",X"eb",X"f3",X"f3",X"0b",X"3c",X"e4",X"0b",X"1b",X"8b",X"39",X"39",X"d1",X"d1",X"d1",X"d1",X"d1",X"57",X"39",X"1f",X"39",X"4a",X"39",X"ae",X"82",X"ae",X"ad",X"1b",X"0b",X"0b",X"ec",X"2e",X"2e",X"d6",X"1b",X"0b",X"2e",X"ea",X"2f",X"2e",X"0b",X"54",X"2e",X"2e",X"75",X"3c",X"25",X"ec",X"4d",X"1b",X"4d",X"2e",X"83",X"0b",X"00",X"00",X"03",X"75",X"03",X"2e",X"75",X"4d",X"ec",X"2e",X"19",X"0b",X"2e",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"27",X"1a",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"00",X"00",X"fb",X"00",X"a4",X"91",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"91",X"f4",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"9e",X"aa",X"92",X"61",X"0b",X"0b",X"0b",X"03",X"03",X"b2",X"03",X"03",X"1a",X"ec",X"2e",X"19",X"19",X"1a",X"1a",X"2f",X"f0",X"f0",X"ed",X"79",X"79",X"61",X"77",X"79",X"54",X"2f",X"f0",X"f0",X"61",X"f0",X"54",X"f0",X"f0",X"28",X"1a",X"03",X"03",X"21",X"03",X"1a",X"03",X"21",X"2e",X"19",X"75",X"75",X"28",X"f0",X"2f",X"79",X"77",X"77",X"79",X"77",X"79",X"f0",X"2f",X"79",X"61",X"79",X"79",X"61",X"77",X"79",X"79",X"75",X"19",X"ec",X"2e",X"2e",X"03",X"1a",X"03",X"cc",X"03",X"1a",X"19",X"28",X"75",X"79",X"61",X"79",X"79",X"61",X"79",X"61",X"79",X"f0",X"f0",X"ed",X"61",X"79",X"77",X"79",X"79",X"79",X"79",X"75",X"19",X"19",X"21",X"2e",X"03",X"1a",X"03",X"b2",X"03",X"0b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"9e",X"aa",X"7c",X"aa",X"61",X"0b",X"0b",X"1b",X"61",X"03",X"b2",X"03",X"b2",X"27",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"71",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"2e",X"0b",X"ed",X"2e",X"0b",X"0b",X"f3",X"6f",X"f3",X"3c",X"0b",X"1a",X"2f",X"0b",X"3c",X"0b",X"65",X"39",X"d1",X"57",X"d1",X"57",X"d1",X"d1",X"39",X"d1",X"39",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"0b",X"3c",X"0b",X"0b",X"2e",X"2e",X"3c",X"0b",X"ec",X"fc",X"0b",X"3c",X"0b",X"ed",X"2e",X"2e",X"fc",X"3c",X"73",X"ec",X"e9",X"00",X"4d",X"2e",X"2e",X"00",X"00",X"00",X"03",X"b2",X"03",X"d6",X"aa",X"60",X"2e",X"2e",X"aa",X"0b",X"2e",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"71",X"19",X"03",X"03",X"75",X"03",X"b2",X"27",X"03",X"1a",X"03",X"b2",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"fb",X"f4",X"fb",X"f4",X"91",X"f4",X"fb",X"f4",X"f4",X"fb",X"f4",X"fb",X"f4",X"4f",X"f4",X"4f",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",X"42",X"6d",X"aa",X"aa",X"84",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"1a",X"03",X"cc",X"19",X"75",X"0d",X"62",X"51",X"cf",X"62",X"62",X"cf",X"62",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"62",X"51",X"62",X"15",X"cf",X"15",X"62",X"62",X"62",X"75",X"75",X"03",X"cc",X"03",X"cc",X"19",X"19",X"75",X"62",X"51",X"62",X"cf",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"cf",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"0d",X"1a",X"03",X"21",X"03",X"21",X"03",X"75",X"75",X"62",X"62",X"51",X"15",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"cf",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"15",X"62",X"75",X"19",X"03",X"cc",X"03",X"1a",X"03",X"19",X"0b",X"3c",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"2f",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"1a",X"03",X"03",X"75",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"2e",X"0b",X"3c",X"2e",X"3c",X"0b",X"4e",X"f3",X"f3",X"0b",X"0b",X"03",X"19",X"2f",X"54",X"1b",X"0b",X"00",X"f3",X"d1",X"d1",X"d1",X"57",X"39",X"1f",X"39",X"4a",X"39",X"ae",X"ae",X"82",X"f3",X"22",X"0b",X"1b",X"0b",X"00",X"d6",X"2e",X"1b",X"0b",X"2e",X"e9",X"00",X"0b",X"00",X"0b",X"ec",X"2e",X"e9",X"1b",X"42",X"ec",X"73",X"1b",X"fc",X"2e",X"1b",X"2e",X"00",X"03",X"19",X"03",X"1a",X"32",X"4d",X"aa",X"2e",X"2e",X"42",X"3c",X"2e",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"71",X"19",X"71",X"03",X"1a",X"03",X"b2",X"19",X"03",X"03",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f4",X"f4",X"fb",X"fb",X"fb",X"f4",X"4f",X"fb",X"91",X"f4",X"4f",X"f4",X"fb",X"f4",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"6d",X"aa",X"9e",X"7c",X"61",X"0b",X"0b",X"1b",X"1a",X"03",X"b2",X"03",X"2e",X"03",X"75",X"15",X"62",X"15",X"f5",X"15",X"f5",X"15",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"62",X"51",X"62",X"75",X"03",X"2e",X"03",X"75",X"62",X"51",X"15",X"62",X"62",X"15",X"51",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"15",X"f5",X"15",X"62",X"51",X"15",X"51",X"62",X"51",X"62",X"15",X"cf",X"19",X"03",X"2e",X"19",X"75",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"1a",X"03",X"2e",X"03",X"b2",X"03",X"0b",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"aa",X"84",X"0b",X"0b",X"0b",X"79",X"03",X"75",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"19",X"03",X"71",X"19",X"71",X"03",X"03",X"19",X"03",X"03",X"1a",X"ec",X"0b",X"1b",X"2e",X"0b",X"3c",X"f3",X"8b",X"46",X"0b",X"3c",X"03",X"b2",X"27",X"ed",X"0b",X"4e",X"0b",X"0b",X"00",X"0b",X"f3",X"d1",X"d1",X"39",X"d1",X"39",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"0b",X"3c",X"0b",X"0b",X"ea",X"2e",X"0b",X"3c",X"2e",X"4d",X"1b",X"1b",X"0b",X"0b",X"0b",X"30",X"4d",X"1b",X"ea",X"2e",X"73",X"3c",X"ea",X"2e",X"1b",X"4d",X"2e",X"03",X"b2",X"03",X"03",X"73",X"e9",X"3c",X"2e",X"ec",X"fc",X"1b",X"2e",X"03",X"03",X"1a",X"03",X"03",X"71",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"fb",X"fb",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"4a",X"f4",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"d8",X"19",X"03",X"03",X"cc",X"1a",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"51",X"cf",X"62",X"62",X"15",X"f5",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"cf",X"62",X"62",X"51",X"75",X"ec",X"75",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"51",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"75",X"ec",X"75",X"15",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"15",X"f5",X"51",X"cf",X"15",X"f5",X"51",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"cf",X"62",X"15",X"cf",X"1a",X"2e",X"03",X"1a",X"03",X"0b",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"9e",X"7c",X"61",X"0b",X"0b",X"1b",X"ed",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"b2",X"19",X"03",X"19",X"b2",X"27",X"19",X"03",X"03",X"1a",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"2e",X"3c",X"0b",X"ec",X"0b",X"1b",X"6f",X"f3",X"f3",X"0b",X"0b",X"1a",X"03",X"b2",X"f0",X"0b",X"39",X"d1",X"0b",X"0b",X"1b",X"0b",X"0b",X"f3",X"d1",X"39",X"4a",X"39",X"ae",X"82",X"ae",X"f3",X"f3",X"1b",X"0b",X"0b",X"0b",X"aa",X"2e",X"3c",X"0b",X"2e",X"d6",X"0b",X"0b",X"00",X"0b",X"00",X"0b",X"0b",X"3c",X"54",X"2e",X"d6",X"0b",X"9e",X"2e",X"0b",X"ea",X"2e",X"1a",X"03",X"19",X"b2",X"fc",X"4d",X"1b",X"d6",X"2e",X"4d",X"1b",X"d6",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"71",X"27",X"19",X"b2",X"03",X"03",X"b2",X"19",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f4",X"f3",X"82",X"70",X"82",X"82",X"70",X"82",X"82",X"70",X"82",X"82",X"82",X"f4",X"f4",X"91",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"9e",X"aa",X"60",X"98",X"0b",X"0b",X"0b",X"19",X"71",X"75",X"ec",X"19",X"15",X"f5",X"51",X"62",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"15",X"f5",X"15",X"51",X"62",X"62",X"62",X"51",X"62",X"cf",X"62",X"15",X"62",X"62",X"51",X"62",X"15",X"cf",X"62",X"51",X"19",X"15",X"51",X"62",X"62",X"51",X"62",X"15",X"f5",X"51",X"62",X"15",X"cf",X"15",X"62",X"62",X"62",X"51",X"62",X"15",X"62",X"cf",X"62",X"15",X"cf",X"15",X"51",X"62",X"62",X"51",X"62",X"62",X"19",X"62",X"51",X"62",X"51",X"62",X"cf",X"15",X"62",X"51",X"cf",X"62",X"15",X"62",X"62",X"15",X"62",X"51",X"62",X"cf",X"62",X"51",X"15",X"cf",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"15",X"75",X"ec",X"03",X"1a",X"1b",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"79",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"03",X"b2",X"19",X"b2",X"03",X"03",X"03",X"75",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"2e",X"1b",X"0b",X"2e",X"0b",X"00",X"f3",X"4e",X"f3",X"0b",X"3c",X"03",X"19",X"03",X"58",X"0b",X"39",X"d1",X"39",X"ae",X"0b",X"3c",X"0b",X"3c",X"0b",X"af",X"39",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"48",X"3c",X"0b",X"1b",X"ed",X"2e",X"0b",X"00",X"2e",X"32",X"1b",X"1b",X"0b",X"00",X"0b",X"0b",X"3c",X"0b",X"ed",X"2e",X"d6",X"1b",X"aa",X"2e",X"3c",X"9e",X"2e",X"03",X"03",X"b2",X"03",X"ea",X"73",X"3c",X"d6",X"2e",X"73",X"3c",X"d6",X"ea",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"03",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"70",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"70",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7f",X"0b",X"cd",X"f0",X"6d",X"f0",X"6d",X"aa",X"7c",X"aa",X"aa",X"33",X"1b",X"0b",X"0b",X"03",X"19",X"03",X"cc",X"1a",X"51",X"15",X"62",X"cf",X"62",X"51",X"cf",X"62",X"51",X"15",X"62",X"62",X"51",X"62",X"62",X"cf",X"15",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"f5",X"62",X"15",X"62",X"28",X"62",X"62",X"15",X"cf",X"62",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"62",X"cf",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"cf",X"15",X"f5",X"62",X"51",X"75",X"15",X"f5",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"cf",X"62",X"62",X"62",X"15",X"62",X"62",X"62",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"75",X"2e",X"19",X"03",X"0b",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"60",X"61",X"0b",X"0b",X"0b",X"2f",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"b2",X"19",X"03",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"2e",X"0b",X"3c",X"2e",X"1b",X"0b",X"65",X"f3",X"f3",X"4e",X"0b",X"03",X"b2",X"27",X"98",X"1b",X"39",X"4a",X"d1",X"57",X"d1",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"00",X"8b",X"ae",X"82",X"f3",X"f3",X"22",X"0b",X"3c",X"0b",X"54",X"2e",X"1b",X"0b",X"2e",X"2e",X"8b",X"4e",X"8b",X"1b",X"0b",X"3c",X"0b",X"0b",X"3c",X"2e",X"2e",X"00",X"f0",X"2e",X"0b",X"2f",X"2e",X"03",X"1a",X"03",X"03",X"1a",X"d6",X"3c",X"e9",X"ec",X"d6",X"1b",X"e9",X"19",X"03",X"19",X"03",X"b2",X"d8",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"b2",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"4f",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",X"9e",X"aa",X"9e",X"7c",X"61",X"0b",X"0b",X"1b",X"19",X"71",X"03",X"e5",X"f0",X"62",X"62",X"62",X"15",X"f5",X"15",X"62",X"62",X"62",X"cf",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"77",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"15",X"f5",X"15",X"f5",X"51",X"62",X"51",X"62",X"62",X"62",X"15",X"51",X"f5",X"79",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"2f",X"2e",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"0d",X"aa",X"98",X"0b",X"0b",X"1b",X"61",X"03",X"75",X"03",X"b2",X"27",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"03",X"b2",X"19",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"2e",X"1b",X"0b",X"2e",X"3c",X"0b",X"f3",X"6f",X"f3",X"6f",X"1b",X"0b",X"03",X"b2",X"2f",X"0b",X"ae",X"57",X"39",X"ff",X"d1",X"3c",X"0b",X"00",X"0b",X"0b",X"3c",X"0b",X"1b",X"0b",X"eb",X"ae",X"f3",X"8b",X"3c",X"0b",X"1b",X"3c",X"2e",X"3c",X"0b",X"2e",X"2e",X"af",X"f3",X"6f",X"f3",X"8b",X"1b",X"0b",X"00",X"0b",X"2e",X"2e",X"0b",X"54",X"2e",X"1b",X"0b",X"2e",X"d6",X"03",X"19",X"b2",X"03",X"d6",X"0b",X"4d",X"2e",X"d6",X"0b",X"4d",X"e9",X"03",X"b2",X"27",X"19",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"6d",X"f0",X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"2e",X"f0",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"62",X"15",X"62",X"51",X"15",X"62",X"62",X"62",X"cf",X"62",X"51",X"62",X"cf",X"15",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"f0",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"f5",X"15",X"cf",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"ed",X"62",X"62",X"15",X"cf",X"62",X"15",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"15",X"62",X"cf",X"62",X"51",X"62",X"62",X"51",X"62",X"2f",X"2e",X"03",X"19",X"0b",X"1b",X"0b",X"3b",X"1a",X"6d",X"3f",X"6d",
    X"9e",X"aa",X"7c",X"aa",X"61",X"0b",X"0b",X"1b",X"2f",X"03",X"b2",X"03",X"19",X"71",X"19",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"19",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"ec",X"0b",X"00",X"2e",X"1b",X"0b",X"4e",X"f3",X"f3",X"ae",X"0b",X"3c",X"19",X"03",X"54",X"00",X"f3",X"fb",X"d1",X"d1",X"d1",X"8b",X"1b",X"0b",X"0b",X"03",X"58",X"54",X"3c",X"0b",X"1b",X"3c",X"f3",X"b8",X"0b",X"0b",X"00",X"2e",X"2e",X"1b",X"0b",X"ec",X"2e",X"6f",X"4e",X"f3",X"f3",X"ae",X"ae",X"8b",X"0b",X"0b",X"ec",X"2e",X"1b",X"2f",X"2e",X"0b",X"3c",X"2f",X"42",X"2e",X"d6",X"03",X"03",X"e5",X"1b",X"42",X"2e",X"ec",X"f0",X"42",X"4d",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"3f",X"f0",X"6d",X"aa",X"12",X"aa",X"2c",X"61",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"2e",X"2f",X"62",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"cf",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"15",X"62",X"62",X"62",X"62",X"cf",X"62",X"62",X"51",X"62",X"51",X"62",X"ed",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"15",X"62",X"cf",X"62",X"62",X"ed",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"cf",X"62",X"62",X"cf",X"62",X"62",X"51",X"62",X"51",X"62",X"cf",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"cf",X"62",X"51",X"62",X"ed",X"2e",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"79",X"03",X"19",X"03",X"b2",X"19",X"03",X"03",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"2e",X"0b",X"0b",X"2e",X"2e",X"00",X"f3",X"4e",X"f3",X"f3",X"ad",X"0b",X"1b",X"03",X"1a",X"1b",X"8b",X"d1",X"39",X"d1",X"57",X"6f",X"3c",X"0b",X"3c",X"19",X"03",X"54",X"1b",X"82",X"8b",X"0b",X"1b",X"0b",X"3c",X"1b",X"2e",X"2e",X"2e",X"00",X"0b",X"2e",X"2e",X"af",X"f3",X"4e",X"f3",X"ae",X"39",X"ae",X"39",X"d1",X"2e",X"2e",X"3c",X"54",X"2e",X"00",X"0b",X"0b",X"54",X"ea",X"42",X"d6",X"2e",X"2e",X"3c",X"ea",X"2e",X"2e",X"54",X"fc",X"f8",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"6d",X"aa",X"aa",X"12",X"98",X"1b",X"0b",X"0b",X"03",X"b2",X"03",X"2e",X"2f",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"62",X"51",X"15",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"51",X"f5",X"15",X"cf",X"62",X"15",X"62",X"62",X"ed",X"62",X"62",X"15",X"cf",X"15",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"62",X"51",X"cf",X"62",X"15",X"cf",X"15",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"f0",X"62",X"62",X"51",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"62",X"62",X"62",X"15",X"62",X"cf",X"15",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"ed",X"2e",X"03",X"19",X"0b",X"0b",X"1b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"84",X"0b",X"0b",X"0b",X"79",X"b2",X"03",X"1a",X"03",X"03",X"19",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"b2",X"d8",X"03",X"1a",X"ec",X"0b",X"1b",X"2e",X"2e",X"46",X"8b",X"f3",X"f3",X"ae",X"f3",X"70",X"0b",X"0b",X"3c",X"0b",X"3c",X"39",X"d1",X"57",X"d1",X"f3",X"1b",X"0b",X"0b",X"03",X"b2",X"f0",X"0b",X"ae",X"f3",X"ae",X"0b",X"3c",X"0b",X"0b",X"2e",X"2e",X"2e",X"1b",X"0b",X"eb",X"2e",X"8b",X"af",X"f3",X"f3",X"ae",X"ae",X"39",X"4a",X"39",X"2e",X"2e",X"1b",X"54",X"2e",X"1b",X"1b",X"0b",X"3c",X"0b",X"1b",X"0b",X"54",X"19",X"1b",X"0b",X"2e",X"2e",X"2f",X"54",X"d6",X"03",X"19",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"b2",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"4a",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"60",X"aa",X"98",X"0b",X"0b",X"1b",X"19",X"03",X"19",X"ec",X"54",X"62",X"15",X"f5",X"51",X"62",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"62",X"cf",X"62",X"15",X"62",X"51",X"15",X"62",X"51",X"62",X"15",X"62",X"15",X"62",X"51",X"62",X"cf",X"62",X"51",X"79",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"51",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"f5",X"51",X"62",X"62",X"51",X"62",X"62",X"cf",X"62",X"51",X"62",X"15",X"62",X"62",X"ed",X"51",X"62",X"62",X"62",X"51",X"62",X"15",X"f5",X"15",X"62",X"51",X"f5",X"cf",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"cf",X"62",X"51",X"15",X"62",X"62",X"51",X"62",X"cf",X"62",X"2f",X"2e",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"9e",X"aa",X"9e",X"7c",X"61",X"0b",X"1b",X"83",X"2f",X"03",X"19",X"03",X"b2",X"19",X"71",X"03",X"19",X"03",X"1a",X"03",X"03",X"75",X"03",X"b2",X"27",X"03",X"1a",X"03",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"19",X"03",X"2e",X"3c",X"0b",X"2e",X"ec",X"8b",X"f3",X"6f",X"f3",X"22",X"ae",X"ae",X"82",X"d1",X"0b",X"1b",X"0b",X"d1",X"d1",X"d1",X"d1",X"ae",X"0b",X"0b",X"00",X"03",X"1a",X"2f",X"0b",X"82",X"ae",X"f3",X"f3",X"0b",X"1b",X"0b",X"3c",X"2e",X"2e",X"3c",X"0b",X"4e",X"8b",X"4e",X"f3",X"6f",X"f3",X"ae",X"39",X"ae",X"39",X"4a",X"2e",X"2e",X"3c",X"ed",X"2e",X"39",X"6f",X"0b",X"1b",X"0b",X"00",X"0b",X"3c",X"0b",X"0b",X"0b",X"d6",X"2e",X"fc",X"2f",X"d6",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"19",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"fb",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"84",X"6d",X"f0",X"6d",X"3f",X"6d",X"42",X"aa",X"9e",X"98",X"0b",X"1b",X"0b",X"03",X"b2",X"03",X"2e",X"54",X"51",X"62",X"62",X"15",X"51",X"62",X"15",X"f5",X"cf",X"62",X"62",X"51",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"f5",X"ed",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"cf",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"15",X"f5",X"51",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"cf",X"62",X"51",X"79",X"62",X"62",X"51",X"cf",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"51",X"f5",X"cf",X"15",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"62",X"cf",X"15",X"62",X"62",X"62",X"51",X"79",X"2e",X"03",X"19",X"0b",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"2f",X"19",X"71",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"b2",X"19",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"2e",X"0b",X"1b",X"2e",X"2e",X"f3",X"4e",X"f3",X"f3",X"ae",X"f3",X"ae",X"ae",X"82",X"39",X"39",X"0b",X"39",X"d1",X"d1",X"57",X"d1",X"0b",X"1b",X"0b",X"00",X"03",X"58",X"0b",X"ae",X"f3",X"ae",X"f3",X"0b",X"3c",X"0b",X"3c",X"2e",X"ec",X"0b",X"1b",X"8b",X"65",X"8b",X"4e",X"f3",X"f3",X"ae",X"ae",X"39",X"d1",X"39",X"2e",X"2e",X"1b",X"0b",X"2e",X"d1",X"39",X"4a",X"ae",X"8b",X"0b",X"1b",X"0b",X"3c",X"0b",X"3c",X"d6",X"2e",X"ea",X"0b",X"2e",X"19",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"4a",X"f4",X"3c",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"3b",X"f0",X"6d",X"f0",X"6d",X"aa",X"2c",X"aa",X"7c",X"61",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"2e",X"2f",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"15",X"51",X"62",X"62",X"15",X"f5",X"15",X"f5",X"15",X"f5",X"62",X"62",X"15",X"62",X"cf",X"62",X"62",X"51",X"62",X"15",X"51",X"f5",X"51",X"79",X"51",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"61",X"51",X"62",X"15",X"f5",X"15",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"f5",X"15",X"62",X"62",X"51",X"62",X"15",X"f5",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"ed",X"2e",X"03",X"b2",X"1b",X"83",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"9e",X"aa",X"60",X"61",X"0b",X"1b",X"0b",X"79",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"ec",X"0b",X"00",X"2e",X"2e",X"8b",X"f3",X"4e",X"f3",X"f3",X"ae",X"82",X"70",X"d1",X"ae",X"39",X"fb",X"57",X"39",X"ff",X"d1",X"d1",X"0b",X"3c",X"0b",X"63",X"00",X"03",X"0b",X"f3",X"ae",X"f3",X"f3",X"0b",X"1b",X"0b",X"0b",X"2e",X"2e",X"f0",X"0b",X"af",X"6f",X"af",X"f3",X"6f",X"f3",X"ae",X"39",X"ae",X"39",X"4a",X"2e",X"2e",X"3c",X"0b",X"2e",X"d1",X"4a",X"39",X"d1",X"82",X"ae",X"8b",X"0b",X"1b",X"0b",X"3c",X"73",X"ec",X"fc",X"1b",X"2e",X"03",X"b2",X"27",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"12",X"aa",X"aa",X"98",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"ec",X"61",X"62",X"51",X"15",X"cf",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"15",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"61",X"62",X"15",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"cf",X"15",X"62",X"51",X"cf",X"15",X"62",X"62",X"62",X"62",X"cf",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"f5",X"62",X"ed",X"62",X"62",X"62",X"51",X"f5",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"15",X"51",X"62",X"51",X"62",X"cf",X"62",X"15",X"62",X"62",X"62",X"15",X"f5",X"62",X"62",X"15",X"51",X"62",X"62",X"ed",X"2e",X"1a",X"03",X"0b",X"3c",X"0b",X"17",X"f0",X"6d",X"f0",X"f0",
    X"aa",X"7c",X"0d",X"aa",X"98",X"0b",X"0b",X"0b",X"79",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"71",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"e5",X"1b",X"0b",X"2e",X"1b",X"0b",X"65",X"f3",X"f3",X"ae",X"f3",X"ae",X"ae",X"ae",X"39",X"39",X"39",X"4a",X"d1",X"d1",X"d1",X"57",X"0b",X"1b",X"0b",X"3c",X"0b",X"00",X"1b",X"8b",X"f3",X"ae",X"f3",X"0b",X"3c",X"0b",X"3c",X"d6",X"2e",X"d6",X"aa",X"98",X"1b",X"8b",X"af",X"f3",X"f3",X"ae",X"82",X"39",X"39",X"d1",X"2e",X"2e",X"1b",X"0b",X"39",X"d1",X"39",X"39",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"0b",X"3c",X"73",X"ec",X"e9",X"3c",X"d6",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"f4",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"6d",X"42",X"60",X"98",X"1b",X"0b",X"1b",X"03",X"b2",X"03",X"2e",X"54",X"62",X"62",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"cf",X"15",X"62",X"62",X"15",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"51",X"2f",X"62",X"51",X"62",X"cf",X"62",X"15",X"62",X"15",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"cf",X"15",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"51",X"79",X"51",X"62",X"15",X"62",X"15",X"62",X"62",X"15",X"cf",X"15",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"62",X"51",X"cf",X"62",X"51",X"62",X"cf",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"2f",X"2e",X"03",X"19",X"0b",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"6d",
    X"9e",X"aa",X"7c",X"aa",X"61",X"0b",X"1b",X"0b",X"ed",X"03",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"d8",X"2e",X"3c",X"0b",X"2e",X"00",X"1b",X"0b",X"00",X"38",X"f3",X"ae",X"ae",X"82",X"39",X"ae",X"39",X"4a",X"57",X"39",X"d1",X"57",X"d1",X"d1",X"39",X"0b",X"1b",X"0b",X"00",X"0b",X"eb",X"ae",X"f3",X"f3",X"0b",X"1b",X"0b",X"0b",X"d6",X"2e",X"00",X"2e",X"d6",X"aa",X"98",X"0b",X"1b",X"f3",X"ae",X"39",X"ae",X"4a",X"39",X"2e",X"2e",X"3c",X"0b",X"d1",X"d1",X"39",X"4a",X"39",X"ae",X"ae",X"ae",X"f3",X"f3",X"0b",X"1b",X"ea",X"2e",X"73",X"3c",X"d6",X"fc",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"75",X"03",X"1a",X"03",X"19",X"b2",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"12",X"aa",X"2c",X"aa",X"23",X"0b",X"0b",X"0b",X"d8",X"1a",X"03",X"2e",X"2f",X"62",X"51",X"62",X"51",X"62",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"cf",X"62",X"62",X"15",X"51",X"62",X"51",X"62",X"cf",X"15",X"62",X"62",X"62",X"ed",X"62",X"62",X"62",X"15",X"62",X"62",X"cf",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"62",X"cf",X"62",X"62",X"51",X"62",X"62",X"53",X"62",X"62",X"51",X"cf",X"62",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"cf",X"62",X"15",X"62",X"54",X"2e",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"f0",
    X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"28",X"03",X"b2",X"03",X"1a",X"03",X"71",X"19",X"71",X"19",X"71",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"19",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"2e",X"0b",X"1b",X"2e",X"0b",X"1a",X"03",X"0b",X"00",X"0b",X"1b",X"38",X"ae",X"ae",X"39",X"39",X"d1",X"39",X"d1",X"57",X"d1",X"d1",X"57",X"d1",X"d1",X"39",X"0b",X"0b",X"1b",X"0b",X"f3",X"ae",X"f3",X"0b",X"3c",X"0b",X"3c",X"42",X"2e",X"00",X"3c",X"3c",X"2e",X"d6",X"aa",X"98",X"0b",X"0b",X"ae",X"39",X"39",X"39",X"2e",X"2e",X"1b",X"0b",X"39",X"d1",X"39",X"d1",X"ae",X"39",X"82",X"f3",X"ae",X"f3",X"0b",X"3c",X"42",X"2e",X"d6",X"1b",X"73",X"4d",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"03",X"1a",X"03",X"b2",X"27",X"03",X"b2",X"03",X"03",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"f0",X"6d",X"f0",X"3f",X"6d",X"42",X"aa",X"9e",X"98",X"0b",X"0b",X"7d",X"19",X"03",X"1a",X"2e",X"2f",X"62",X"62",X"15",X"62",X"51",X"15",X"62",X"62",X"cf",X"15",X"f5",X"51",X"62",X"15",X"cf",X"62",X"62",X"51",X"62",X"15",X"cf",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"cf",X"15",X"62",X"53",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"15",X"f5",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"51",X"15",X"cf",X"15",X"51",X"62",X"77",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"cf",X"62",X"15",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"62",X"62",X"15",X"62",X"cf",X"62",X"2f",X"2e",X"03",X"19",X"1b",X"0b",X"1b",X"17",X"3f",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"84",X"0b",X"0b",X"0b",X"77",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"75",X"03",X"03",X"b2",X"19",X"71",X"27",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"2e",X"2f",X"0b",X"2e",X"1b",X"03",X"0b",X"0b",X"1b",X"0b",X"00",X"0b",X"00",X"eb",X"ae",X"39",X"fb",X"d1",X"d1",X"d1",X"d1",X"57",X"d1",X"39",X"d1",X"39",X"39",X"4a",X"0b",X"0b",X"ae",X"f3",X"f3",X"8b",X"1b",X"0b",X"0b",X"ea",X"2e",X"00",X"00",X"e9",X"00",X"00",X"2e",X"d6",X"aa",X"0b",X"1b",X"4e",X"39",X"fb",X"d1",X"2e",X"2e",X"1b",X"d1",X"39",X"fb",X"39",X"39",X"ae",X"ae",X"ae",X"f3",X"f3",X"48",X"3c",X"0b",X"32",X"d6",X"0b",X"4d",X"e9",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"6d",X"aa",X"aa",X"2c",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"b2",X"03",X"2e",X"ed",X"62",X"51",X"62",X"cf",X"62",X"62",X"51",X"62",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"f0",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"62",X"62",X"cf",X"15",X"62",X"62",X"62",X"51",X"15",X"62",X"62",X"cf",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"ed",X"62",X"62",X"62",X"51",X"62",X"cf",X"62",X"15",X"f5",X"51",X"62",X"62",X"62",X"15",X"62",X"cf",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"79",X"2e",X"03",X"b2",X"0b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"9e",X"7c",X"61",X"0b",X"0b",X"1b",X"2f",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"71",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"e5",X"54",X"1b",X"d6",X"1b",X"0b",X"3c",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"3c",X"eb",X"39",X"39",X"d1",X"57",X"d1",X"d1",X"d1",X"d1",X"d1",X"4a",X"39",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"4e",X"0b",X"3c",X"0b",X"9e",X"2e",X"00",X"00",X"2e",X"2e",X"d6",X"aa",X"54",X"1b",X"3c",X"0b",X"0b",X"0b",X"39",X"d1",X"d1",X"2e",X"d1",X"39",X"d1",X"39",X"39",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"22",X"1b",X"0b",X"e9",X"ec",X"0b",X"fc",X"4d",X"19",X"71",X"19",X"71",X"27",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"4a",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"6d",X"f0",X"aa",X"12",X"aa",X"92",X"61",X"0b",X"0b",X"0b",X"19",X"03",X"19",X"2e",X"2f",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"cf",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"ed",X"51",X"62",X"15",X"62",X"51",X"15",X"cf",X"62",X"62",X"51",X"62",X"51",X"cf",X"62",X"51",X"62",X"62",X"62",X"51",X"15",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"f0",X"51",X"62",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"51",X"f5",X"62",X"15",X"62",X"cf",X"62",X"51",X"62",X"cf",X"62",X"15",X"62",X"62",X"62",X"15",X"62",X"53",X"2e",X"1a",X"03",X"0b",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"0b",X"83",X"28",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"03",X"1a",X"03",X"19",X"b2",X"19",X"71",X"19",X"71",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"2e",X"aa",X"0b",X"32",X"0b",X"1b",X"6f",X"f3",X"f3",X"ae",X"f3",X"8b",X"0b",X"00",X"0b",X"0b",X"0b",X"3c",X"eb",X"d1",X"57",X"d1",X"57",X"39",X"d1",X"39",X"39",X"d1",X"82",X"ae",X"ae",X"f3",X"f3",X"f3",X"0b",X"1b",X"0b",X"aa",X"2e",X"2e",X"d6",X"aa",X"54",X"1b",X"0b",X"3c",X"0b",X"8b",X"39",X"ae",X"39",X"4a",X"d1",X"39",X"d1",X"ff",X"d1",X"d1",X"39",X"fb",X"39",X"ae",X"82",X"ae",X"f3",X"f3",X"f3",X"0b",X"0b",X"4d",X"2e",X"2f",X"42",X"d6",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"03",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"3f",X"f0",X"6d",X"aa",X"2c",X"aa",X"aa",X"98",X"1b",X"0b",X"1b",X"03",X"b2",X"03",X"2e",X"2f",X"62",X"51",X"62",X"15",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"cf",X"15",X"62",X"51",X"62",X"cf",X"15",X"62",X"15",X"51",X"62",X"15",X"62",X"ed",X"62",X"62",X"cf",X"62",X"62",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"15",X"62",X"15",X"cf",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"cf",X"15",X"62",X"62",X"62",X"15",X"62",X"62",X"ed",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"cf",X"15",X"62",X"15",X"51",X"62",X"51",X"62",X"15",X"62",X"62",X"15",X"62",X"62",X"cf",X"62",X"51",X"62",X"62",X"ed",X"2e",X"03",X"03",X"0b",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"9e",X"aa",X"60",X"61",X"0b",X"1b",X"0b",X"2f",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"03",X"19",X"03",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"2e",X"aa",X"0b",X"73",X"3c",X"4e",X"f3",X"f3",X"f3",X"f3",X"ae",X"82",X"b7",X"8b",X"1b",X"0b",X"3c",X"0b",X"0b",X"0b",X"0b",X"d1",X"d1",X"d1",X"d1",X"39",X"4a",X"82",X"39",X"ae",X"f3",X"ae",X"f3",X"4e",X"0b",X"00",X"0b",X"aa",X"2e",X"3c",X"0b",X"1b",X"0b",X"3c",X"1b",X"6f",X"f3",X"ae",X"82",X"39",X"39",X"d1",X"39",X"d1",X"ff",X"d1",X"39",X"d1",X"39",X"39",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"8b",X"3c",X"1b",X"fc",X"2e",X"f0",X"54",X"d6",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"03",X"b2",X"19",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"4a",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"54",X"f0",X"6d",X"3f",X"aa",X"12",X"aa",X"6d",X"23",X"0b",X"0b",X"0b",X"03",X"1a",X"03",X"2e",X"54",X"62",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"cf",X"62",X"15",X"62",X"15",X"62",X"51",X"62",X"15",X"f5",X"51",X"62",X"cf",X"62",X"62",X"62",X"cf",X"62",X"2f",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"62",X"cf",X"15",X"51",X"62",X"cf",X"15",X"61",X"51",X"62",X"62",X"cf",X"62",X"62",X"62",X"15",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"79",X"2e",X"03",X"1a",X"e4",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"0d",X"aa",X"98",X"0b",X"0b",X"0b",X"79",X"03",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"75",X"03",X"b2",X"19",X"b2",X"27",X"75",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"cc",X"aa",X"0b",X"4d",X"2e",X"f3",X"f3",X"22",X"f3",X"ae",X"f3",X"ae",X"ae",X"82",X"8b",X"3c",X"0b",X"0b",X"3c",X"3c",X"e4",X"1b",X"0b",X"39",X"d1",X"39",X"d1",X"39",X"ae",X"82",X"ae",X"f3",X"f3",X"f3",X"0b",X"0b",X"0b",X"ed",X"2e",X"0b",X"00",X"0b",X"8b",X"af",X"6f",X"f3",X"f3",X"ae",X"39",X"ae",X"39",X"39",X"1f",X"39",X"d1",X"d1",X"d1",X"d1",X"39",X"4a",X"39",X"ae",X"ae",X"82",X"f3",X"0b",X"3c",X"0b",X"0b",X"42",X"2e",X"42",X"2f",X"2e",X"74",X"33",X"03",X"1a",X"03",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"53",X"6d",X"3f",X"6d",X"f0",X"2c",X"aa",X"92",X"aa",X"84",X"0b",X"0b",X"1b",X"19",X"03",X"1a",X"2e",X"2f",X"62",X"51",X"62",X"62",X"15",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"62",X"cf",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"77",X"62",X"62",X"15",X"62",X"15",X"51",X"62",X"62",X"cf",X"62",X"62",X"62",X"cf",X"62",X"62",X"62",X"62",X"cf",X"15",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"ed",X"62",X"62",X"51",X"62",X"15",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"cf",X"15",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"cf",X"15",X"f5",X"51",X"61",X"2e",X"03",X"19",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",
    X"9e",X"aa",X"7c",X"aa",X"61",X"0b",X"0b",X"1b",X"ed",X"03",X"19",X"b2",X"03",X"1a",X"03",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"2e",X"fc",X"0b",X"fc",X"2e",X"f3",X"6f",X"f3",X"46",X"f3",X"ae",X"82",X"70",X"d1",X"ae",X"8b",X"1b",X"0b",X"0b",X"0b",X"1a",X"00",X"0b",X"3c",X"0b",X"4a",X"39",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"6f",X"3c",X"1b",X"0b",X"2f",X"2e",X"1b",X"0b",X"4e",X"eb",X"8b",X"f3",X"4e",X"f3",X"ae",X"ae",X"39",X"4a",X"d1",X"39",X"d1",X"ff",X"d1",X"39",X"d1",X"39",X"d1",X"82",X"39",X"ae",X"0b",X"0b",X"00",X"0b",X"0b",X"3c",X"ea",X"ec",X"fc",X"1b",X"2e",X"00",X"74",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"75",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"12",X"aa",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"b2",X"03",X"2e",X"2f",X"62",X"62",X"62",X"51",X"62",X"cf",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"15",X"f5",X"62",X"15",X"f5",X"ed",X"62",X"51",X"62",X"62",X"cf",X"62",X"15",X"51",X"62",X"15",X"62",X"51",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"62",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"ed",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"cf",X"62",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"ed",X"2e",X"03",X"b2",X"1b",X"0b",X"1b",X"17",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"2f",X"03",X"b2",X"03",X"03",X"19",X"71",X"19",X"b2",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"71",X"19",X"b2",X"27",X"19",X"03",X"2e",X"ea",X"0b",X"42",X"2e",X"af",X"f3",X"f3",X"f3",X"ae",X"f3",X"ae",X"ae",X"82",X"39",X"4a",X"0b",X"3c",X"0b",X"00",X"03",X"0b",X"0b",X"0b",X"00",X"0b",X"3c",X"0b",X"ae",X"82",X"ae",X"f3",X"f3",X"f3",X"0b",X"0b",X"3c",X"98",X"2e",X"0b",X"3c",X"8b",X"4e",X"8b",X"4e",X"f3",X"f3",X"ae",X"39",X"ae",X"39",X"39",X"d1",X"39",X"d1",X"ff",X"d1",X"d1",X"4a",X"39",X"4a",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"3c",X"2e",X"2e",X"e9",X"3c",X"d6",X"23",X"00",X"84",X"03",X"b2",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"19",X"71",X"19",X"71",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"91",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"79",X"6d",X"f0",X"6d",X"aa",X"60",X"aa",X"7c",X"33",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"2e",X"2f",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"cf",X"15",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"15",X"51",X"62",X"15",X"cf",X"15",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"53",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"15",X"51",X"62",X"62",X"cf",X"15",X"51",X"62",X"15",X"62",X"15",X"62",X"61",X"62",X"15",X"51",X"62",X"cf",X"15",X"62",X"62",X"15",X"cf",X"15",X"62",X"15",X"f5",X"51",X"62",X"62",X"51",X"62",X"15",X"62",X"cf",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"f0",X"2e",X"1a",X"03",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"84",X"0b",X"0b",X"1b",X"79",X"03",X"1a",X"03",X"19",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"03",X"19",X"71",X"19",X"03",X"19",X"03",X"71",X"19",X"03",X"71",X"19",X"03",X"03",X"b2",X"03",X"1a",X"ec",X"42",X"1b",X"aa",X"2e",X"2e",X"4e",X"f3",X"f3",X"f3",X"ae",X"ae",X"70",X"d1",X"ae",X"39",X"eb",X"0b",X"1b",X"0b",X"0b",X"1b",X"f3",X"d1",X"f3",X"8b",X"1b",X"0b",X"3c",X"0b",X"f3",X"ae",X"f3",X"6f",X"3c",X"0b",X"3c",X"0b",X"2e",X"f0",X"0b",X"6f",X"af",X"8b",X"f3",X"4e",X"f3",X"ae",X"ae",X"39",X"39",X"fb",X"39",X"d1",X"57",X"d1",X"39",X"d1",X"39",X"1b",X"0b",X"0b",X"3c",X"0b",X"0b",X"1b",X"2f",X"42",X"2e",X"2e",X"2e",X"4d",X"1b",X"32",X"42",X"00",X"74",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"b2",X"27",X"03",X"b2",X"03",X"19",X"03",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"f0",X"3f",X"6d",X"aa",X"aa",X"12",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"b2",X"03",X"2e",X"ed",X"62",X"62",X"15",X"51",X"f5",X"62",X"15",X"62",X"62",X"cf",X"15",X"f5",X"51",X"a1",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"62",X"cf",X"15",X"62",X"62",X"cf",X"15",X"62",X"51",X"62",X"2f",X"62",X"51",X"62",X"62",X"51",X"15",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"cf",X"62",X"62",X"51",X"79",X"51",X"62",X"62",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"cf",X"15",X"f5",X"51",X"15",X"62",X"51",X"62",X"ed",X"2e",X"03",X"19",X"0b",X"1b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"9e",X"7c",X"61",X"0b",X"0b",X"0b",X"2f",X"19",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"75",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"e5",X"bc",X"0b",X"aa",X"2e",X"2e",X"f3",X"f3",X"22",X"ae",X"f3",X"82",X"ae",X"82",X"39",X"d1",X"39",X"6f",X"00",X"0b",X"0b",X"f3",X"d1",X"d1",X"39",X"4a",X"39",X"48",X"1b",X"0b",X"0b",X"f3",X"22",X"f3",X"1b",X"0b",X"00",X"0b",X"ec",X"aa",X"0b",X"af",X"8b",X"4e",X"8b",X"f3",X"f3",X"ae",X"39",X"ae",X"39",X"39",X"d1",X"d1",X"d1",X"d1",X"57",X"0b",X"00",X"0b",X"0b",X"3c",X"0b",X"3c",X"2f",X"42",X"2e",X"2e",X"2e",X"ec",X"2e",X"d6",X"0b",X"e9",X"d8",X"0a",X"00",X"23",X"03",X"b2",X"19",X"b2",X"03",X"19",X"03",X"b2",X"19",X"03",X"19",X"71",X"19",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"2c",X"aa",X"aa",X"23",X"0b",X"0b",X"0b",X"19",X"03",X"19",X"2e",X"2f",X"f5",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"15",X"f5",X"51",X"8e",X"51",X"62",X"62",X"62",X"15",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"15",X"f5",X"51",X"62",X"15",X"f5",X"58",X"62",X"62",X"15",X"62",X"62",X"62",X"cf",X"15",X"62",X"00",X"62",X"62",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"15",X"61",X"62",X"62",X"51",X"15",X"62",X"62",X"15",X"f5",X"62",X"51",X"f5",X"51",X"62",X"62",X"cf",X"15",X"f5",X"51",X"a1",X"62",X"62",X"51",X"62",X"62",X"62",X"15",X"62",X"62",X"62",X"cf",X"62",X"2f",X"2e",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"6d",X"3f",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"28",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"d6",X"73",X"1b",X"9e",X"2e",X"2e",X"4e",X"f3",X"f3",X"f3",X"ae",X"ae",X"ae",X"39",X"ae",X"39",X"d1",X"d1",X"0b",X"1b",X"b8",X"57",X"d1",X"39",X"ff",X"39",X"4a",X"ae",X"82",X"8b",X"3c",X"0b",X"f3",X"f3",X"0b",X"0b",X"0b",X"0b",X"2e",X"4d",X"1b",X"0b",X"4e",X"8b",X"f3",X"6f",X"f3",X"ae",X"ae",X"39",X"d1",X"4a",X"39",X"d1",X"57",X"d1",X"1b",X"0b",X"1b",X"0b",X"3c",X"0b",X"0b",X"2e",X"2e",X"32",X"74",X"00",X"2e",X"2e",X"2e",X"d6",X"3c",X"4d",X"e9",X"61",X"00",X"74",X"1a",X"03",X"03",X"03",X"19",X"b2",X"27",X"19",X"03",X"03",X"b2",X"d8",X"19",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"12",X"aa",X"60",X"98",X"0b",X"1b",X"0b",X"03",X"19",X"71",X"2e",X"2f",X"62",X"62",X"51",X"62",X"62",X"cf",X"62",X"62",X"62",X"62",X"51",X"18",X"8e",X"f5",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"15",X"f5",X"cf",X"62",X"ed",X"62",X"62",X"51",X"cf",X"15",X"51",X"62",X"51",X"1b",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"15",X"62",X"51",X"62",X"ed",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"15",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"51",X"f5",X"8e",X"a1",X"62",X"62",X"15",X"51",X"62",X"cf",X"62",X"51",X"62",X"15",X"62",X"53",X"2e",X"03",X"19",X"0b",X"0b",X"1b",X"3b",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"9e",X"aa",X"60",X"61",X"0b",X"0b",X"0b",X"79",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"d6",X"4d",X"1b",X"2f",X"2e",X"2e",X"f3",X"f3",X"6f",X"0b",X"00",X"0b",X"65",X"ae",X"39",X"39",X"4a",X"39",X"f3",X"0b",X"ff",X"d1",X"d1",X"57",X"87",X"39",X"ae",X"39",X"ae",X"82",X"0b",X"1b",X"0b",X"3c",X"0b",X"3c",X"1b",X"3c",X"2e",X"2e",X"3c",X"0b",X"eb",X"8b",X"4e",X"f3",X"f3",X"ae",X"39",X"ae",X"39",X"39",X"d1",X"39",X"d1",X"d1",X"d1",X"0b",X"0b",X"1b",X"0b",X"3c",X"0b",X"ed",X"54",X"fc",X"2e",X"2e",X"2e",X"ec",X"2e",X"2e",X"1b",X"42",X"73",X"ba",X"00",X"74",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"4f",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"cd",X"6d",X"f0",X"6d",X"f0",X"60",X"aa",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"19",X"71",X"19",X"2e",X"2f",X"62",X"15",X"cf",X"62",X"51",X"62",X"51",X"62",X"51",X"51",X"de",X"8e",X"8e",X"a1",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"f5",X"51",X"62",X"51",X"62",X"15",X"62",X"ed",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"62",X"3c",X"62",X"00",X"23",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"62",X"62",X"cf",X"15",X"51",X"62",X"cf",X"62",X"62",X"ed",X"62",X"62",X"62",X"cf",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"51",X"62",X"15",X"51",X"62",X"51",X"8e",X"18",X"51",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"ed",X"2e",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"7c",X"0d",X"aa",X"98",X"0b",X"1b",X"0b",X"77",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"71",X"fc",X"d6",X"0b",X"54",X"2e",X"2e",X"4e",X"f3",X"3c",X"1b",X"0b",X"2d",X"1b",X"f3",X"ae",X"39",X"d1",X"d1",X"39",X"f3",X"d1",X"d1",X"57",X"4a",X"57",X"39",X"39",X"ae",X"82",X"b7",X"f3",X"6f",X"00",X"0b",X"0b",X"0b",X"2e",X"2e",X"33",X"2e",X"1b",X"0b",X"8b",X"af",X"f3",X"4e",X"f3",X"ae",X"ae",X"39",X"fb",X"39",X"d1",X"d1",X"d1",X"57",X"39",X"1f",X"39",X"39",X"0b",X"1b",X"0b",X"00",X"0b",X"0b",X"54",X"2f",X"42",X"2e",X"2e",X"2e",X"3c",X"42",X"d6",X"74",X"74",X"00",X"33",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"75",X"03",X"1a",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"aa",X"2c",X"12",X"98",X"1b",X"0b",X"0b",X"27",X"75",X"03",X"cc",X"54",X"51",X"62",X"62",X"15",X"62",X"15",X"f5",X"62",X"51",X"18",X"8e",X"8e",X"18",X"a1",X"34",X"0f",X"0f",X"f5",X"41",X"a9",X"41",X"41",X"41",X"41",X"41",X"41",X"62",X"62",X"62",X"51",X"62",X"ed",X"62",X"15",X"f5",X"51",X"62",X"51",X"62",X"51",X"62",X"3c",X"4b",X"00",X"12",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"51",X"62",X"15",X"f5",X"62",X"62",X"62",X"51",X"62",X"53",X"62",X"51",X"15",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"a1",X"18",X"8e",X"de",X"51",X"62",X"51",X"62",X"15",X"62",X"15",X"62",X"62",X"51",X"f0",X"2e",X"03",X"19",X"0b",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"7c",X"aa",X"61",X"0b",X"0b",X"0b",X"79",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"75",X"03",X"b2",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"ea",X"d6",X"00",X"2f",X"2e",X"2e",X"f3",X"f3",X"0b",X"0b",X"2d",X"a5",X"63",X"1b",X"39",X"4a",X"39",X"39",X"8a",X"d1",X"57",X"d1",X"d1",X"ff",X"39",X"fb",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"0b",X"1b",X"0b",X"00",X"2e",X"b6",X"1b",X"2e",X"3c",X"0b",X"eb",X"4e",X"8b",X"f3",X"f3",X"ae",X"39",X"ae",X"39",X"39",X"d1",X"d1",X"d1",X"57",X"d1",X"39",X"39",X"fb",X"39",X"39",X"0b",X"0b",X"0b",X"1b",X"3c",X"0b",X"0b",X"ed",X"54",X"ea",X"3c",X"1b",X"d6",X"00",X"00",X"00",X"74",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"03",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"92",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"b2",X"03",X"03",X"2e",X"2f",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"18",X"8e",X"8e",X"8e",X"8e",X"18",X"24",X"18",X"24",X"18",X"18",X"5b",X"18",X"24",X"18",X"18",X"b1",X"41",X"62",X"51",X"15",X"62",X"62",X"ed",X"51",X"62",X"62",X"15",X"62",X"62",X"15",X"62",X"00",X"12",X"00",X"00",X"4b",X"12",X"00",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"15",X"51",X"f0",X"62",X"62",X"f5",X"51",X"62",X"41",X"41",X"41",X"41",X"41",X"41",X"a9",X"f5",X"a9",X"34",X"0f",X"51",X"0f",X"8e",X"8e",X"8e",X"18",X"a1",X"62",X"51",X"62",X"51",X"cf",X"62",X"51",X"62",X"ed",X"2e",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"1b",X"61",X"b2",X"03",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"19",X"03",X"19",X"b2",X"27",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"2e",X"0b",X"0b",X"2e",X"2e",X"4e",X"f3",X"0b",X"1b",X"0b",X"0b",X"33",X"0b",X"eb",X"39",X"d1",X"4a",X"39",X"d1",X"ff",X"d1",X"57",X"39",X"d1",X"39",X"39",X"ae",X"82",X"ae",X"f3",X"f3",X"6f",X"3c",X"0b",X"0b",X"3c",X"2e",X"1b",X"2e",X"1b",X"0b",X"4e",X"8b",X"f3",X"4e",X"f3",X"ae",X"82",X"39",X"39",X"fb",X"39",X"d1",X"d1",X"d1",X"39",X"d1",X"d1",X"39",X"fb",X"ae",X"39",X"ae",X"ae",X"0b",X"0b",X"1b",X"0b",X"3c",X"0b",X"0b",X"0b",X"0b",X"ea",X"d6",X"4c",X"00",X"84",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"19",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"3f",X"6d",X"aa",X"aa",X"9e",X"98",X"0b",X"0b",X"3c",X"19",X"03",X"1a",X"ec",X"54",X"62",X"51",X"62",X"62",X"62",X"51",X"51",X"18",X"8e",X"8e",X"8e",X"8e",X"8e",X"18",X"8e",X"18",X"24",X"18",X"5b",X"18",X"30",X"18",X"30",X"5b",X"8e",X"41",X"51",X"62",X"62",X"cf",X"62",X"ed",X"62",X"62",X"51",X"62",X"51",X"62",X"cf",X"62",X"00",X"23",X"2e",X"4b",X"12",X"23",X"00",X"23",X"23",X"74",X"00",X"00",X"00",X"00",X"62",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"53",X"62",X"51",X"15",X"62",X"f5",X"41",X"8e",X"8e",X"18",X"18",X"24",X"18",X"24",X"18",X"9a",X"18",X"24",X"8e",X"8e",X"8e",X"8e",X"8e",X"18",X"a1",X"62",X"62",X"62",X"62",X"15",X"62",X"62",X"2f",X"2e",X"03",X"19",X"0b",X"0b",X"3c",X"17",X"6d",X"f0",X"6d",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"84",X"0b",X"0b",X"0b",X"2f",X"03",X"03",X"1a",X"03",X"19",X"71",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"2e",X"1b",X"0b",X"65",X"2e",X"f3",X"f3",X"4e",X"0b",X"0b",X"1b",X"0b",X"3c",X"0b",X"ae",X"39",X"39",X"d1",X"39",X"d1",X"d1",X"d1",X"d1",X"39",X"fb",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"f3",X"1b",X"0b",X"1b",X"0b",X"2e",X"7f",X"33",X"2e",X"3c",X"0b",X"65",X"8b",X"f3",X"f3",X"ae",X"39",X"ae",X"39",X"39",X"d1",X"d1",X"d1",X"57",X"d1",X"39",X"4a",X"39",X"39",X"39",X"ae",X"ae",X"70",X"f3",X"ae",X"0b",X"1b",X"0b",X"3c",X"0b",X"3c",X"0b",X"ed",X"d6",X"ed",X"74",X"00",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"12",X"aa",X"7c",X"61",X"0b",X"1b",X"0b",X"03",X"b2",X"03",X"2e",X"ed",X"62",X"62",X"15",X"62",X"cf",X"3a",X"8f",X"8e",X"41",X"8e",X"8e",X"8e",X"18",X"8e",X"18",X"24",X"18",X"5b",X"18",X"5b",X"8f",X"c7",X"8f",X"c7",X"18",X"41",X"62",X"62",X"51",X"62",X"15",X"61",X"62",X"51",X"62",X"cf",X"62",X"15",X"62",X"51",X"3c",X"00",X"12",X"12",X"23",X"00",X"23",X"ba",X"23",X"23",X"23",X"00",X"00",X"00",X"62",X"51",X"62",X"cf",X"62",X"15",X"0f",X"62",X"62",X"2f",X"62",X"62",X"62",X"cf",X"15",X"41",X"8e",X"c7",X"5b",X"18",X"30",X"18",X"24",X"18",X"24",X"18",X"18",X"8e",X"18",X"8e",X"8e",X"8e",X"8e",X"18",X"51",X"51",X"62",X"51",X"62",X"cf",X"62",X"ed",X"2e",X"b2",X"03",X"0b",X"1b",X"0b",X"33",X"f0",X"6d",X"3f",X"f0",
    X"9e",X"aa",X"9e",X"7c",X"61",X"0b",X"1b",X"0b",X"79",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"19",X"03",X"75",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"2e",X"0b",X"3c",X"4e",X"8b",X"4e",X"f3",X"f3",X"46",X"ae",X"f3",X"8b",X"0b",X"1b",X"39",X"4a",X"39",X"d1",X"d1",X"57",X"f3",X"0b",X"3c",X"0b",X"39",X"39",X"ae",X"ae",X"82",X"82",X"f3",X"22",X"48",X"3c",X"0b",X"3c",X"0b",X"2e",X"33",X"ba",X"2e",X"3c",X"1b",X"0b",X"eb",X"f3",X"ae",X"ae",X"39",X"4a",X"d1",X"39",X"d1",X"ff",X"d1",X"39",X"8a",X"39",X"39",X"fb",X"ae",X"39",X"ae",X"82",X"ae",X"f3",X"f3",X"8b",X"f3",X"1b",X"0b",X"0b",X"3c",X"54",X"2e",X"00",X"f8",X"00",X"03",X"75",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"79",X"6d",X"f0",X"6d",X"9e",X"aa",X"2c",X"aa",X"84",X"0b",X"0b",X"0b",X"19",X"03",X"19",X"2e",X"2f",X"62",X"51",X"62",X"62",X"51",X"51",X"41",X"8e",X"be",X"8e",X"8e",X"8e",X"8e",X"f9",X"8e",X"18",X"18",X"24",X"18",X"30",X"18",X"30",X"18",X"30",X"8e",X"41",X"62",X"51",X"62",X"62",X"62",X"ed",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"3c",X"23",X"00",X"00",X"00",X"12",X"12",X"12",X"23",X"23",X"ba",X"00",X"00",X"3c",X"62",X"15",X"62",X"51",X"62",X"cf",X"62",X"15",X"51",X"54",X"51",X"62",X"51",X"62",X"62",X"41",X"8e",X"c7",X"30",X"8f",X"c7",X"30",X"18",X"5b",X"18",X"45",X"18",X"24",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"18",X"51",X"62",X"62",X"51",X"62",X"15",X"61",X"2e",X"03",X"19",X"0b",X"0b",X"0b",X"3b",X"3f",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"0b",X"0b",X"ed",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"d8",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"cc",X"3c",X"0b",X"8b",X"af",X"f3",X"6f",X"f3",X"f3",X"f3",X"ae",X"ae",X"ae",X"0b",X"ae",X"39",X"4a",X"d1",X"39",X"d1",X"0b",X"1b",X"0b",X"2e",X"0b",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"f3",X"f3",X"0b",X"1b",X"0b",X"00",X"2e",X"33",X"74",X"63",X"2e",X"2e",X"1b",X"3c",X"0b",X"ae",X"39",X"ae",X"39",X"39",X"1f",X"39",X"d1",X"d1",X"d1",X"39",X"39",X"4a",X"39",X"39",X"ae",X"82",X"ae",X"f3",X"ae",X"f3",X"f3",X"4e",X"0b",X"0b",X"00",X"0b",X"1b",X"2e",X"00",X"f8",X"00",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"12",X"aa",X"98",X"56",X"0b",X"1b",X"03",X"b2",X"03",X"2e",X"98",X"62",X"62",X"51",X"15",X"62",X"62",X"51",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"18",X"18",X"24",X"18",X"24",X"9a",X"24",X"c7",X"8f",X"30",X"8f",X"b1",X"41",X"62",X"62",X"51",X"62",X"51",X"79",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"00",X"23",X"23",X"12",X"12",X"12",X"12",X"12",X"12",X"23",X"23",X"ba",X"00",X"3c",X"51",X"62",X"51",X"62",X"15",X"62",X"15",X"cf",X"62",X"2f",X"62",X"62",X"15",X"51",X"62",X"41",X"8e",X"5b",X"30",X"18",X"8f",X"18",X"8f",X"18",X"18",X"24",X"18",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"be",X"41",X"51",X"62",X"51",X"62",X"62",X"62",X"77",X"2e",X"03",X"b2",X"5d",X"0b",X"0b",X"98",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"60",X"61",X"0b",X"3c",X"0b",X"79",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"19",X"b2",X"19",X"03",X"19",X"71",X"19",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"2e",X"1b",X"0b",X"65",X"48",X"4e",X"f3",X"f3",X"f3",X"ae",X"f3",X"ae",X"70",X"ae",X"39",X"d1",X"39",X"39",X"8a",X"d1",X"0b",X"00",X"e5",X"c7",X"ee",X"0b",X"82",X"ae",X"82",X"82",X"f3",X"22",X"af",X"0b",X"0b",X"3c",X"0b",X"0b",X"2e",X"23",X"b6",X"3b",X"6a",X"2e",X"2e",X"1b",X"0b",X"0b",X"39",X"4a",X"39",X"39",X"d1",X"ff",X"d1",X"d1",X"d1",X"39",X"d1",X"39",X"ae",X"39",X"ae",X"ae",X"ae",X"f3",X"f3",X"4e",X"f3",X"0b",X"1b",X"0b",X"0b",X"3c",X"2e",X"2f",X"74",X"00",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"3b",X"6d",X"3f",X"6d",X"f0",X"7c",X"aa",X"9e",X"aa",X"98",X"1b",X"0b",X"0b",X"19",X"03",X"1a",X"ec",X"2f",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"51",X"41",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"18",X"8e",X"18",X"18",X"45",X"18",X"8e",X"41",X"62",X"51",X"62",X"62",X"15",X"98",X"62",X"62",X"62",X"15",X"62",X"51",X"62",X"cf",X"7a",X"23",X"23",X"12",X"2e",X"12",X"12",X"12",X"12",X"23",X"23",X"23",X"3c",X"3c",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"ed",X"62",X"51",X"62",X"62",X"62",X"41",X"8e",X"21",X"c7",X"5b",X"c7",X"24",X"9a",X"18",X"24",X"18",X"8e",X"18",X"8e",X"8e",X"8e",X"8e",X"8e",X"41",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"ed",X"2e",X"19",X"03",X"0b",X"0b",X"1b",X"3b",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"0d",X"aa",X"98",X"0b",X"83",X"0b",X"2f",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"2e",X"00",X"0b",X"1b",X"38",X"f3",X"f3",X"22",X"f3",X"f3",X"ae",X"82",X"ae",X"39",X"ae",X"39",X"4a",X"d1",X"39",X"d1",X"0b",X"1b",X"0b",X"2d",X"2d",X"4c",X"0b",X"82",X"ae",X"ae",X"f3",X"f3",X"f3",X"8b",X"3c",X"0b",X"0b",X"3c",X"2e",X"33",X"b6",X"c6",X"00",X"b6",X"b6",X"2e",X"ec",X"3c",X"0b",X"0b",X"3c",X"d1",X"39",X"d1",X"57",X"d1",X"39",X"4a",X"39",X"fb",X"39",X"ae",X"ae",X"70",X"f3",X"ae",X"f3",X"f3",X"8b",X"1b",X"3c",X"0b",X"3c",X"0b",X"2e",X"b1",X"00",X"74",X"03",X"b2",X"27",X"1a",X"03",X"03",X"b2",X"27",X"19",X"b2",X"03",X"1a",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"60",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"03",X"b2",X"03",X"2e",X"54",X"62",X"15",X"62",X"cf",X"62",X"62",X"15",X"62",X"51",X"41",X"8e",X"8e",X"18",X"a1",X"51",X"a1",X"f5",X"0f",X"0f",X"f5",X"f5",X"34",X"f5",X"41",X"41",X"41",X"62",X"15",X"62",X"cf",X"62",X"ed",X"62",X"51",X"62",X"cf",X"62",X"15",X"51",X"62",X"51",X"3c",X"23",X"12",X"12",X"12",X"12",X"12",X"12",X"23",X"23",X"23",X"3c",X"51",X"62",X"51",X"cf",X"15",X"51",X"62",X"62",X"51",X"62",X"77",X"62",X"62",X"62",X"cf",X"15",X"41",X"8e",X"18",X"24",X"18",X"8e",X"18",X"8e",X"8e",X"8e",X"18",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"51",X"51",X"62",X"15",X"cf",X"62",X"51",X"62",X"77",X"2e",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"9e",X"aa",X"7c",X"aa",X"61",X"0b",X"0b",X"1b",X"79",X"03",X"75",X"03",X"b2",X"d8",X"03",X"75",X"03",X"19",X"03",X"71",X"19",X"03",X"19",X"03",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"75",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"2e",X"1b",X"0b",X"00",X"0b",X"eb",X"f3",X"f3",X"ae",X"82",X"ae",X"ae",X"82",X"39",X"39",X"d1",X"39",X"1f",X"57",X"f3",X"0b",X"1b",X"0b",X"3c",X"4c",X"0b",X"0b",X"82",X"f3",X"ae",X"f3",X"4e",X"f3",X"0b",X"3c",X"0b",X"0b",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"1b",X"00",X"0b",X"3c",X"0b",X"eb",X"d1",X"39",X"d1",X"d1",X"39",X"39",X"ae",X"39",X"ae",X"ae",X"ae",X"f3",X"f3",X"4e",X"f3",X"0b",X"0b",X"3c",X"0b",X"3c",X"2e",X"00",X"00",X"74",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"19",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"4f",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"7c",X"9e",X"98",X"0b",X"1b",X"0b",X"19",X"03",X"19",X"2e",X"2f",X"f5",X"51",X"62",X"62",X"15",X"cf",X"62",X"51",X"62",X"51",X"41",X"8e",X"8e",X"51",X"62",X"62",X"15",X"cf",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"62",X"51",X"62",X"51",X"15",X"51",X"79",X"62",X"62",X"15",X"51",X"62",X"62",X"15",X"62",X"62",X"3c",X"23",X"23",X"12",X"12",X"12",X"12",X"23",X"23",X"23",X"3c",X"3c",X"62",X"62",X"15",X"62",X"62",X"62",X"cf",X"15",X"f5",X"51",X"79",X"51",X"62",X"51",X"62",X"62",X"f5",X"f5",X"f5",X"41",X"f5",X"41",X"0f",X"f5",X"f5",X"a1",X"51",X"a1",X"f5",X"8e",X"8e",X"8e",X"41",X"a1",X"51",X"62",X"51",X"62",X"62",X"62",X"15",X"f5",X"ed",X"2e",X"03",X"19",X"0b",X"1b",X"0b",X"33",X"f0",X"6d",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"2f",X"03",X"b2",X"03",X"19",X"b2",X"19",X"71",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"ec",X"2e",X"1b",X"0b",X"0b",X"0b",X"3c",X"4e",X"82",X"ae",X"39",X"ae",X"4a",X"39",X"d1",X"39",X"d1",X"d1",X"57",X"d1",X"6f",X"1b",X"0b",X"3c",X"1b",X"0b",X"ae",X"f3",X"f3",X"f3",X"4e",X"0b",X"1b",X"0b",X"00",X"2e",X"1b",X"0b",X"00",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"00",X"0b",X"0b",X"0b",X"3c",X"0b",X"00",X"0b",X"0b",X"eb",X"39",X"4a",X"39",X"ae",X"82",X"ae",X"f3",X"ae",X"f3",X"f3",X"6f",X"00",X"0b",X"0b",X"0b",X"00",X"2e",X"84",X"00",X"33",X"03",X"03",X"19",X"03",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"f4",X"f4",X"3c",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"53",X"6d",X"f0",X"3f",X"6d",X"6d",X"aa",X"9e",X"aa",X"98",X"0b",X"0b",X"0b",X"d8",X"b2",X"03",X"2e",X"2f",X"f5",X"15",X"f5",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"41",X"8e",X"0f",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"15",X"cf",X"62",X"62",X"62",X"62",X"62",X"61",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"3c",X"3c",X"23",X"23",X"23",X"23",X"23",X"3c",X"3c",X"3c",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"f5",X"61",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"f5",X"51",X"8e",X"8e",X"8e",X"51",X"62",X"15",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"79",X"2e",X"03",X"b2",X"1b",X"0b",X"0b",X"53",X"6d",X"f0",X"3f",X"54",
    X"aa",X"7c",X"aa",X"aa",X"84",X"0b",X"1b",X"0b",X"77",X"03",X"19",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"03",X"1a",X"2e",X"00",X"0b",X"00",X"0b",X"0b",X"3c",X"f3",X"ae",X"39",X"39",X"d1",X"39",X"d1",X"57",X"d1",X"d1",X"d1",X"ff",X"39",X"fb",X"6f",X"0b",X"e4",X"f3",X"ae",X"f3",X"4e",X"f3",X"6f",X"3c",X"3c",X"0b",X"0b",X"3c",X"0b",X"0b",X"00",X"0b",X"0b",X"3c",X"0b",X"0b",X"0b",X"0b",X"3c",X"3c",X"0b",X"3c",X"0b",X"0b",X"00",X"0b",X"0b",X"3c",X"0b",X"39",X"ae",X"82",X"ae",X"f3",X"22",X"8b",X"f3",X"1b",X"0b",X"00",X"0b",X"0b",X"2e",X"00",X"74",X"03",X"19",X"b2",X"19",X"71",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"aa",X"7c",X"aa",X"61",X"0b",X"0b",X"1b",X"19",X"03",X"1a",X"2e",X"2f",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"51",X"41",X"51",X"62",X"62",X"51",X"62",X"51",X"cf",X"15",X"62",X"51",X"62",X"51",X"62",X"51",X"15",X"62",X"51",X"62",X"2f",X"62",X"62",X"62",X"62",X"cf",X"15",X"f5",X"62",X"51",X"15",X"62",X"62",X"3c",X"00",X"00",X"3c",X"3c",X"3c",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"15",X"f5",X"51",X"62",X"51",X"2f",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"15",X"cf",X"15",X"62",X"62",X"51",X"62",X"62",X"51",X"51",X"18",X"8e",X"51",X"51",X"62",X"cf",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"ed",X"2e",X"03",X"19",X"0b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"6d",
    X"9e",X"aa",X"9e",X"7c",X"61",X"0b",X"0b",X"83",X"2f",X"03",X"b2",X"03",X"19",X"03",X"19",X"b2",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"19",X"2e",X"2e",X"3c",X"0b",X"1b",X"0b",X"0b",X"00",X"0b",X"0b",X"0b",X"0b",X"f3",X"4a",X"d1",X"d1",X"d1",X"d1",X"57",X"d1",X"39",X"d1",X"39",X"39",X"ae",X"ae",X"82",X"f3",X"f3",X"f3",X"6f",X"af",X"0b",X"0b",X"0b",X"00",X"0b",X"0b",X"1b",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"1b",X"3c",X"0b",X"0b",X"0b",X"3c",X"0b",X"1b",X"0b",X"00",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"00",X"82",X"f3",X"f3",X"4e",X"0b",X"3c",X"0b",X"3c",X"1b",X"2e",X"00",X"ba",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"0d",X"12",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"03",X"b2",X"03",X"2e",X"ed",X"62",X"51",X"62",X"15",X"cf",X"62",X"15",X"62",X"cf",X"62",X"62",X"cf",X"0a",X"0f",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"cf",X"62",X"62",X"62",X"62",X"62",X"62",X"cf",X"62",X"51",X"79",X"51",X"62",X"15",X"51",X"62",X"62",X"15",X"cf",X"62",X"62",X"62",X"51",X"62",X"cf",X"62",X"15",X"62",X"51",X"f5",X"51",X"62",X"cf",X"15",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"62",X"ed",X"62",X"62",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"51",X"41",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"cf",X"15",X"62",X"62",X"62",X"ed",X"2e",X"03",X"b2",X"1b",X"0b",X"3c",X"98",X"f0",X"6d",X"f0",X"3f",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"ed",X"03",X"75",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"03",X"b2",X"19",X"71",X"19",X"03",X"b2",X"2e",X"1b",X"0b",X"1b",X"0b",X"00",X"0b",X"1b",X"0b",X"0b",X"1b",X"1b",X"0b",X"3c",X"0b",X"f3",X"d1",X"d1",X"ff",X"d1",X"d1",X"d1",X"d1",X"39",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"4e",X"f3",X"8b",X"0b",X"3c",X"0b",X"1b",X"38",X"af",X"8b",X"4e",X"f3",X"4e",X"48",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"3c",X"0b",X"0b",X"00",X"0b",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"0b",X"0b",X"3c",X"2e",X"84",X"00",X"b0",X"1a",X"03",X"19",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"3b",X"6d",X"f0",X"6d",X"f0",X"7c",X"aa",X"aa",X"aa",X"98",X"0b",X"0b",X"3c",X"19",X"03",X"19",X"2e",X"2f",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"51",X"cf",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"61",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"cf",X"62",X"15",X"f5",X"15",X"f5",X"51",X"62",X"62",X"15",X"62",X"62",X"62",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"cf",X"62",X"2f",X"62",X"51",X"62",X"62",X"51",X"cf",X"15",X"62",X"f5",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"51",X"51",X"62",X"15",X"62",X"15",X"62",X"51",X"15",X"62",X"62",X"51",X"62",X"ed",X"2e",X"03",X"19",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"79",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"0b",X"0b",X"00",X"0b",X"eb",X"8b",X"f3",X"4e",X"f3",X"ae",X"f3",X"6f",X"0b",X"1b",X"0b",X"00",X"0b",X"3c",X"f3",X"d1",X"57",X"39",X"d1",X"39",X"4a",X"82",X"ae",X"82",X"82",X"f3",X"f3",X"8b",X"4e",X"3c",X"0b",X"3c",X"0b",X"4e",X"8b",X"4e",X"f3",X"6f",X"f3",X"f3",X"ae",X"ae",X"ae",X"82",X"f3",X"6f",X"1b",X"0b",X"0b",X"1b",X"0b",X"00",X"0b",X"00",X"0b",X"00",X"0b",X"3c",X"0b",X"1b",X"0b",X"00",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"2e",X"ba",X"03",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"2c",X"aa",X"12",X"98",X"0b",X"1b",X"0b",X"d8",X"b2",X"03",X"2e",X"f0",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"cf",X"62",X"15",X"62",X"62",X"62",X"62",X"51",X"77",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"15",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"62",X"62",X"62",X"51",X"77",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"15",X"62",X"62",X"62",X"15",X"cf",X"15",X"62",X"15",X"62",X"62",X"62",X"62",X"51",X"62",X"cf",X"62",X"62",X"62",X"62",X"cf",X"15",X"62",X"61",X"2e",X"03",X"b2",X"5d",X"0b",X"0b",X"33",X"6d",X"3f",X"6d",X"f0",
    X"aa",X"7c",X"0d",X"aa",X"84",X"0b",X"0b",X"1b",X"2f",X"03",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"2e",X"2e",X"3c",X"1b",X"6f",X"af",X"8b",X"4e",X"8b",X"f3",X"f3",X"f3",X"ae",X"82",X"70",X"d1",X"f3",X"0b",X"0b",X"1b",X"0b",X"3c",X"b8",X"d1",X"39",X"d1",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"4e",X"f3",X"6f",X"1b",X"0b",X"0b",X"00",X"8b",X"af",X"8b",X"4e",X"f3",X"f3",X"ae",X"f3",X"70",X"d1",X"ae",X"39",X"39",X"1f",X"39",X"ae",X"f3",X"8b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"00",X"0b",X"3c",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"2e",X"33",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"19",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"f0",X"6d",X"6d",X"f0",X"60",X"aa",X"9e",X"aa",X"98",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"ec",X"54",X"15",X"f5",X"51",X"cf",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"cf",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"cf",X"15",X"51",X"f5",X"77",X"62",X"62",X"15",X"cf",X"62",X"15",X"62",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"cf",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"ed",X"f5",X"51",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"cf",X"62",X"51",X"62",X"cf",X"15",X"62",X"62",X"62",X"51",X"62",X"51",X"f5",X"51",X"62",X"51",X"79",X"2e",X"19",X"03",X"0b",X"0b",X"1b",X"17",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"7c",X"aa",X"98",X"0b",X"0b",X"83",X"2f",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"03",X"1a",X"ec",X"0b",X"0b",X"8b",X"af",X"8b",X"4e",X"8b",X"f3",X"6f",X"f3",X"ae",X"f3",X"ae",X"ae",X"82",X"39",X"39",X"fb",X"f3",X"0b",X"1b",X"1b",X"0b",X"3c",X"65",X"39",X"ae",X"ae",X"ae",X"f3",X"f3",X"f3",X"8b",X"af",X"0b",X"3c",X"0b",X"3c",X"6f",X"af",X"6f",X"f3",X"8b",X"f3",X"f3",X"ae",X"ae",X"82",X"39",X"d1",X"d1",X"39",X"57",X"d1",X"57",X"4a",X"57",X"39",X"4a",X"ae",X"8b",X"8b",X"1b",X"0b",X"0b",X"1b",X"0b",X"3c",X"0b",X"00",X"0b",X"3c",X"0b",X"2e",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"b2",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"70",X"3c",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"f3",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"53",X"6d",X"f0",X"3f",X"54",X"42",X"aa",X"7c",X"aa",X"74",X"1b",X"0b",X"3c",X"03",X"b2",X"03",X"2e",X"98",X"62",X"62",X"15",X"f5",X"51",X"62",X"62",X"cf",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"62",X"cf",X"15",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"61",X"62",X"51",X"62",X"62",X"15",X"cf",X"62",X"62",X"51",X"62",X"cf",X"62",X"62",X"62",X"15",X"f5",X"15",X"cf",X"15",X"62",X"62",X"15",X"f5",X"51",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"61",X"15",X"62",X"62",X"62",X"cf",X"15",X"62",X"62",X"cf",X"15",X"62",X"62",X"f5",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"62",X"15",X"62",X"15",X"f5",X"ed",X"2e",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"9e",X"98",X"1b",X"0b",X"1b",X"2f",X"19",X"03",X"1a",X"03",X"03",X"b2",X"d8",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"03",X"b2",X"19",X"03",X"2e",X"0b",X"00",X"eb",X"8b",X"4e",X"8b",X"af",X"4e",X"f3",X"f3",X"f3",X"ae",X"ae",X"70",X"d1",X"ae",X"39",X"39",X"4a",X"d1",X"f3",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"65",X"f3",X"ae",X"f3",X"4e",X"f3",X"4e",X"0b",X"0b",X"0b",X"3c",X"8b",X"eb",X"8b",X"af",X"f3",X"22",X"ae",X"f3",X"ae",X"39",X"ae",X"39",X"39",X"1f",X"d1",X"d1",X"d1",X"ff",X"39",X"4a",X"39",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"22",X"48",X"f3",X"0b",X"0b",X"00",X"0b",X"0b",X"2e",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"82",X"82",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"82",X"70",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"6d",X"aa",X"9e",X"aa",X"98",X"0b",X"0b",X"0b",X"19",X"03",X"19",X"ec",X"2f",X"62",X"51",X"62",X"15",X"f5",X"51",X"62",X"62",X"15",X"cf",X"15",X"62",X"15",X"f5",X"62",X"51",X"62",X"62",X"62",X"62",X"cf",X"62",X"62",X"51",X"62",X"15",X"f5",X"51",X"62",X"51",X"62",X"ed",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"cf",X"62",X"15",X"62",X"62",X"62",X"62",X"cf",X"62",X"62",X"15",X"53",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"cf",X"15",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"f5",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"2f",X"2e",X"03",X"19",X"0b",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"33",X"0b",X"0b",X"0b",X"77",X"03",X"71",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"b2",X"19",X"03",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"2e",X"1b",X"0b",X"4e",X"8b",X"af",X"4e",X"8b",X"f3",X"8b",X"f3",X"ae",X"f3",X"ae",X"82",X"ae",X"39",X"39",X"fb",X"57",X"39",X"d1",X"d1",X"ff",X"f3",X"0b",X"1b",X"3c",X"0b",X"0b",X"65",X"f3",X"f3",X"6f",X"8b",X"00",X"0b",X"3c",X"0b",X"4e",X"8b",X"4e",X"f3",X"6f",X"f3",X"f3",X"ae",X"82",X"ae",X"39",X"4a",X"57",X"39",X"d1",X"ff",X"d1",X"39",X"d1",X"39",X"d1",X"39",X"ae",X"82",X"ae",X"f3",X"f3",X"f3",X"f3",X"4e",X"0b",X"1b",X"0b",X"0b",X"00",X"3c",X"2e",X"03",X"b2",X"03",X"75",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"b2",X"03",X"1a",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f4",X"82",X"82",X"82",X"82",X"82",X"82",X"70",X"82",X"82",X"82",X"82",X"82",X"4a",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"7c",X"aa",X"60",X"98",X"1b",X"0b",X"1b",X"03",X"b2",X"03",X"2e",X"54",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"cf",X"62",X"51",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"62",X"ed",X"62",X"62",X"15",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"15",X"f5",X"51",X"62",X"15",X"f5",X"51",X"cf",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"61",X"62",X"62",X"62",X"15",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"cf",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"79",X"2e",X"b2",X"03",X"0b",X"0b",X"0b",X"3b",X"3f",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"9e",X"7c",X"61",X"0b",X"1b",X"0b",X"f0",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"b2",X"03",X"75",X"03",X"03",X"b2",X"19",X"71",X"19",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"2e",X"3c",X"0b",X"8b",X"af",X"6f",X"8b",X"4e",X"8b",X"46",X"f3",X"f3",X"ae",X"82",X"ae",X"39",X"ae",X"39",X"39",X"39",X"d1",X"ff",X"d1",X"39",X"1f",X"39",X"fb",X"8b",X"0b",X"1b",X"0b",X"0b",X"00",X"0b",X"eb",X"1b",X"0b",X"0b",X"3c",X"0b",X"eb",X"8b",X"af",X"f3",X"f3",X"ae",X"f3",X"ae",X"39",X"ae",X"39",X"d1",X"d1",X"d1",X"57",X"d1",X"ff",X"39",X"4a",X"39",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"46",X"8b",X"f3",X"4e",X"0b",X"3c",X"0b",X"0b",X"0b",X"2e",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"fb",X"f4",X"4f",X"fb",X"f4",X"fb",X"f4",X"91",X"f4",X"4f",X"f4",X"fb",X"f4",X"91",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"3b",X"6d",X"f0",X"6d",X"3f",X"aa",X"9e",X"aa",X"aa",X"84",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"2e",X"2f",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"cf",X"62",X"15",X"f5",X"51",X"62",X"15",X"62",X"cf",X"15",X"62",X"62",X"62",X"62",X"51",X"62",X"ed",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"cf",X"15",X"62",X"62",X"cf",X"15",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"79",X"51",X"62",X"51",X"62",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"cf",X"15",X"51",X"cf",X"15",X"62",X"cf",X"62",X"62",X"51",X"62",X"51",X"cf",X"15",X"62",X"62",X"51",X"62",X"61",X"2e",X"03",X"19",X"0b",X"1b",X"0b",X"53",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"2f",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"06",X"19",X"03",X"03",X"cc",X"2e",X"2e",X"2e",X"03",X"19",X"71",X"03",X"1a",X"03",X"75",X"03",X"b2",X"2e",X"0b",X"1b",X"3c",X"eb",X"8b",X"af",X"eb",X"f3",X"8b",X"22",X"ae",X"f3",X"b7",X"82",X"ae",X"39",X"d1",X"4a",X"d1",X"39",X"57",X"d1",X"57",X"39",X"39",X"39",X"39",X"ae",X"ae",X"8b",X"1b",X"0b",X"0b",X"00",X"0b",X"0b",X"3c",X"0b",X"3c",X"8b",X"4e",X"f3",X"6f",X"f3",X"f3",X"ae",X"82",X"ae",X"39",X"39",X"d1",X"39",X"57",X"d1",X"d1",X"39",X"d1",X"d1",X"39",X"fb",X"ae",X"82",X"ae",X"f3",X"f3",X"f3",X"f3",X"6f",X"af",X"0b",X"0b",X"3c",X"0b",X"3c",X"2e",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"19",X"b2",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f4",X"fb",X"f4",X"f4",X"fb",X"f4",X"fb",X"f4",X"f4",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"00",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"7c",X"9e",X"7c",X"33",X"1b",X"0b",X"1b",X"03",X"b2",X"03",X"2e",X"ed",X"62",X"62",X"15",X"cf",X"62",X"62",X"62",X"62",X"15",X"62",X"62",X"15",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"cf",X"62",X"51",X"62",X"51",X"cf",X"62",X"51",X"62",X"62",X"51",X"f0",X"62",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"cf",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"15",X"f5",X"51",X"62",X"62",X"62",X"51",X"62",X"15",X"98",X"62",X"15",X"62",X"cf",X"62",X"15",X"cf",X"62",X"15",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"51",X"15",X"62",X"15",X"62",X"62",X"62",X"cf",X"15",X"62",X"62",X"ed",X"2e",X"03",X"b2",X"1b",X"0b",X"0b",X"98",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"79",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"03",X"cc",X"2e",X"1b",X"0b",X"3c",X"0b",X"2e",X"2e",X"03",X"1a",X"03",X"03",X"71",X"19",X"03",X"75",X"ec",X"0b",X"0b",X"4e",X"8b",X"4e",X"8b",X"4e",X"f3",X"f3",X"f3",X"ae",X"82",X"ae",X"39",X"ae",X"39",X"39",X"d1",X"d1",X"d1",X"d1",X"39",X"1f",X"d1",X"4a",X"ae",X"39",X"ae",X"f3",X"ae",X"6f",X"1b",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"4e",X"8b",X"4e",X"f3",X"46",X"ae",X"f3",X"ae",X"39",X"ae",X"39",X"4a",X"d1",X"d1",X"d1",X"ff",X"d1",X"39",X"4a",X"39",X"39",X"39",X"ae",X"82",X"ae",X"f3",X"f3",X"4e",X"f3",X"8b",X"1b",X"3c",X"0b",X"3c",X"0b",X"21",X"03",X"b2",X"19",X"03",X"b2",X"27",X"03",X"03",X"75",X"03",X"b2",X"03",X"b2",X"03",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f4",X"fb",X"f4",X"fb",X"91",X"f4",X"4f",X"fb",X"fb",X"fb",X"91",X"f4",X"fb",X"f4",X"fb",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"f0",X"6d",X"f0",X"6d",X"12",X"aa",X"aa",X"aa",X"98",X"0b",X"0b",X"0b",X"19",X"03",X"19",X"2e",X"2f",X"62",X"51",X"62",X"15",X"62",X"cf",X"15",X"51",X"cf",X"62",X"51",X"62",X"62",X"15",X"f5",X"62",X"62",X"15",X"51",X"f5",X"51",X"62",X"62",X"62",X"62",X"62",X"15",X"62",X"cf",X"15",X"62",X"ed",X"62",X"51",X"f5",X"51",X"62",X"62",X"15",X"62",X"62",X"62",X"62",X"15",X"51",X"62",X"51",X"cf",X"62",X"62",X"cf",X"62",X"15",X"62",X"51",X"62",X"15",X"62",X"cf",X"15",X"62",X"cf",X"62",X"ed",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"cf",X"62",X"62",X"51",X"62",X"62",X"51",X"15",X"62",X"62",X"62",X"62",X"cf",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"79",X"2e",X"03",X"19",X"0b",X"0b",X"0b",X"3b",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"84",X"0b",X"1b",X"0b",X"ed",X"03",X"b2",X"19",X"03",X"19",X"71",X"19",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"2e",X"3c",X"0b",X"54",X"f0",X"6d",X"f0",X"0b",X"0b",X"2e",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"2e",X"0b",X"00",X"0b",X"eb",X"8b",X"af",X"f3",X"6f",X"f3",X"ae",X"f3",X"ae",X"ae",X"82",X"39",X"fb",X"39",X"d1",X"39",X"ff",X"d1",X"d1",X"39",X"39",X"39",X"39",X"ae",X"82",X"b7",X"f3",X"f3",X"f3",X"8b",X"1b",X"0b",X"0b",X"0b",X"3c",X"0b",X"eb",X"f3",X"8b",X"f3",X"f3",X"ae",X"82",X"b7",X"8b",X"1b",X"0b",X"1b",X"0b",X"f3",X"d1",X"d1",X"ff",X"39",X"39",X"fb",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"f3",X"6f",X"af",X"0b",X"0b",X"0b",X"0b",X"2e",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"19",X"71",X"27",X"19",X"03",X"19",X"03",X"00",X"00",X"f4",X"3c",X"8f",X"4f",X"f4",X"91",X"f4",X"fb",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"fb",X"f4",X"91",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",X"aa",X"6d",X"aa",X"12",X"98",X"0b",X"1b",X"0b",X"03",X"b2",X"03",X"2e",X"2f",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"15",X"cf",X"62",X"62",X"15",X"62",X"62",X"15",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"f0",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"62",X"15",X"51",X"62",X"62",X"cf",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"15",X"61",X"51",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"f5",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"f5",X"51",X"62",X"ed",X"2e",X"03",X"b2",X"5d",X"0b",X"0b",X"33",X"6d",X"3f",X"6d",X"f0",
    X"9e",X"aa",X"7c",X"9e",X"98",X"0b",X"0b",X"0b",X"79",X"03",X"75",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"27",X"19",X"03",X"2e",X"0b",X"2f",X"98",X"3f",X"6d",X"f0",X"6d",X"f0",X"3f",X"3c",X"2e",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"e5",X"1b",X"0b",X"0b",X"4e",X"8b",X"4e",X"f3",X"f3",X"d7",X"ae",X"82",X"70",X"d1",X"ae",X"39",X"39",X"fb",X"d1",X"d1",X"57",X"d1",X"d1",X"39",X"4a",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"4e",X"8b",X"00",X"0b",X"3c",X"0b",X"00",X"0b",X"00",X"4e",X"f3",X"f3",X"22",X"82",X"ae",X"82",X"ae",X"39",X"0b",X"3c",X"0b",X"0b",X"0b",X"00",X"39",X"d1",X"d1",X"39",X"39",X"ae",X"ae",X"82",X"f3",X"f3",X"6f",X"f3",X"65",X"0b",X"1b",X"0b",X"1b",X"2e",X"03",X"1a",X"03",X"03",X"b2",X"19",X"71",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"00",X"00",X"fb",X"00",X"a4",X"4f",X"f4",X"fb",X"f4",X"fb",X"f4",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"f4",X"fb",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"12",X"aa",X"7c",X"aa",X"84",X"0b",X"0b",X"0b",X"d8",X"1a",X"03",X"2e",X"54",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"cf",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"15",X"f5",X"62",X"51",X"62",X"62",X"ed",X"62",X"62",X"62",X"cf",X"62",X"51",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"51",X"15",X"f5",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"ed",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"15",X"cf",X"62",X"62",X"62",X"15",X"62",X"62",X"15",X"62",X"15",X"51",X"62",X"62",X"15",X"f5",X"ed",X"2e",X"19",X"03",X"0b",X"0b",X"1b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"1b",X"83",X"2f",X"03",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"03",X"b2",X"19",X"b2",X"03",X"2e",X"00",X"2f",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"6d",X"98",X"1b",X"2e",X"03",X"2e",X"2e",X"2e",X"2e",X"2e",X"03",X"2e",X"1b",X"0b",X"3c",X"38",X"f3",X"4e",X"f3",X"f3",X"f3",X"ae",X"ae",X"ae",X"39",X"39",X"4a",X"57",X"39",X"d1",X"d1",X"d1",X"39",X"d1",X"39",X"4a",X"ae",X"ae",X"82",X"f3",X"f3",X"f3",X"4e",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"0b",X"0b",X"eb",X"f3",X"f3",X"ae",X"f3",X"ae",X"39",X"ae",X"39",X"6f",X"1b",X"0b",X"3c",X"0b",X"d1",X"39",X"4a",X"39",X"ae",X"39",X"6f",X"3c",X"0b",X"0b",X"3c",X"1b",X"0b",X"0b",X"3c",X"cc",X"2e",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"19",X"03",X"19",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"f4",X"fb",X"fb",X"00",X"00",X"82",X"82",X"82",X"82",X"82",X"82",X"70",X"3c",X"00",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"aa",X"9e",X"aa",X"98",X"0b",X"1b",X"0b",X"19",X"03",X"1a",X"ec",X"ed",X"62",X"62",X"15",X"cf",X"15",X"51",X"62",X"15",X"f5",X"62",X"15",X"62",X"cf",X"15",X"62",X"51",X"62",X"51",X"62",X"cf",X"15",X"62",X"cf",X"15",X"62",X"cf",X"15",X"62",X"15",X"cf",X"62",X"2f",X"51",X"62",X"51",X"62",X"15",X"f5",X"15",X"62",X"62",X"cf",X"15",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"cf",X"15",X"f5",X"51",X"62",X"62",X"62",X"ed",X"62",X"51",X"62",X"cf",X"15",X"62",X"cf",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"51",X"cf",X"62",X"51",X"62",X"62",X"cf",X"62",X"62",X"62",X"51",X"62",X"62",X"2f",X"2e",X"03",X"b2",X"1b",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"7c",X"aa",X"60",X"ba",X"0b",X"0b",X"1b",X"2f",X"27",X"19",X"03",X"03",X"b2",X"03",X"03",X"19",X"03",X"03",X"03",X"e5",X"1b",X"54",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"6d",X"f0",X"aa",X"aa",X"54",X"2e",X"2e",X"0b",X"0b",X"1b",X"3c",X"0b",X"2e",X"2e",X"ec",X"0b",X"1b",X"0b",X"65",X"f3",X"f3",X"f3",X"ae",X"f3",X"82",X"39",X"ae",X"39",X"d1",X"39",X"d1",X"ff",X"d1",X"39",X"d1",X"4a",X"39",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"4e",X"8b",X"1b",X"3c",X"0b",X"3c",X"0b",X"1b",X"0b",X"3c",X"0b",X"b8",X"f3",X"f3",X"ae",X"82",X"ae",X"39",X"39",X"8a",X"39",X"0b",X"1b",X"0b",X"4a",X"57",X"39",X"4a",X"39",X"ae",X"8b",X"3c",X"0b",X"3c",X"0b",X"0b",X"0b",X"ec",X"2e",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"03",X"03",X"b2",X"00",X"00",X"fb",X"00",X"a4",X"4f",X"fb",X"f4",X"f4",X"3c",X"a4",X"82",X"3c",X"3c",X"3c",X"3c",X"3c",X"82",X"82",X"3c",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"cd",X"6d",X"f0",X"6d",X"f0",X"60",X"aa",X"7c",X"aa",X"61",X"0b",X"0b",X"1b",X"03",X"b2",X"03",X"2e",X"54",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"cf",X"15",X"51",X"f5",X"51",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"53",X"62",X"62",X"15",X"f5",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"cf",X"15",X"51",X"62",X"15",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"ed",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"cf",X"15",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"62",X"f5",X"15",X"f5",X"51",X"62",X"51",X"62",X"cf",X"15",X"62",X"cf",X"15",X"98",X"2e",X"03",X"19",X"0b",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"9e",X"aa",X"98",X"0b",X"1b",X"0b",X"79",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"ec",X"0b",X"54",X"3f",X"f0",X"6d",X"6d",X"f0",X"6d",X"f0",X"60",X"aa",X"92",X"aa",X"0b",X"00",X"54",X"aa",X"a7",X"68",X"d6",X"d6",X"3c",X"42",X"2e",X"2e",X"3c",X"0b",X"0b",X"4e",X"f3",X"f3",X"f3",X"ae",X"ae",X"ae",X"39",X"39",X"4a",X"d1",X"39",X"d1",X"ff",X"d1",X"d1",X"39",X"39",X"39",X"ae",X"82",X"ae",X"f3",X"f3",X"f3",X"6f",X"8b",X"3c",X"0b",X"0b",X"3c",X"0b",X"ec",X"0b",X"3c",X"0b",X"f3",X"ae",X"f3",X"ae",X"39",X"ae",X"39",X"39",X"d1",X"d1",X"57",X"0b",X"ff",X"39",X"4a",X"39",X"ae",X"39",X"ae",X"0b",X"1b",X"0b",X"2e",X"ec",X"2e",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"19",X"03",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"19",X"00",X"00",X"f4",X"3c",X"8f",X"4f",X"f4",X"3c",X"00",X"82",X"82",X"3c",X"a4",X"8f",X"a4",X"8f",X"a4",X"3c",X"82",X"70",X"3c",X"f4",X"3c",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"19",X"03",X"19",X"ec",X"2f",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"15",X"62",X"62",X"62",X"62",X"51",X"62",X"51",X"15",X"51",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"ed",X"62",X"51",X"62",X"51",X"15",X"62",X"62",X"51",X"62",X"15",X"51",X"62",X"62",X"62",X"cf",X"62",X"62",X"15",X"62",X"62",X"15",X"f5",X"62",X"51",X"62",X"62",X"51",X"cf",X"15",X"62",X"62",X"ed",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"15",X"51",X"62",X"62",X"15",X"62",X"62",X"15",X"51",X"62",X"51",X"62",X"62",X"ed",X"2e",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"2f",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"2e",X"0b",X"2f",X"6d",X"f0",X"6d",X"3f",X"54",X"aa",X"1b",X"0b",X"aa",X"aa",X"aa",X"6d",X"a7",X"a7",X"a7",X"0c",X"0c",X"d6",X"d6",X"2e",X"1b",X"0b",X"2e",X"00",X"0b",X"0b",X"7d",X"0b",X"f3",X"46",X"ae",X"f3",X"ae",X"70",X"ae",X"39",X"d1",X"39",X"1f",X"57",X"d1",X"39",X"d1",X"39",X"fb",X"ae",X"39",X"ae",X"f3",X"ae",X"82",X"6f",X"f3",X"4e",X"0b",X"0b",X"3c",X"0b",X"0b",X"2e",X"2e",X"1b",X"0b",X"1b",X"b8",X"ae",X"82",X"ae",X"39",X"fb",X"d1",X"39",X"ff",X"d1",X"d1",X"39",X"d1",X"d1",X"39",X"39",X"ae",X"ae",X"0b",X"3c",X"0b",X"2e",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"b2",X"03",X"03",X"00",X"00",X"fb",X"00",X"a4",X"4f",X"3c",X"8f",X"00",X"82",X"3c",X"a4",X"8f",X"a4",X"8f",X"a4",X"a4",X"8f",X"00",X"82",X"3c",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"b2",X"03",X"2e",X"98",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"cf",X"51",X"15",X"cf",X"15",X"62",X"62",X"62",X"62",X"62",X"51",X"15",X"62",X"51",X"62",X"51",X"15",X"cf",X"15",X"62",X"ed",X"62",X"62",X"15",X"f5",X"cf",X"62",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"cf",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"ed",X"62",X"62",X"62",X"15",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"cf",X"15",X"51",X"cf",X"62",X"15",X"f5",X"51",X"cf",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"51",X"79",X"2e",X"03",X"19",X"0b",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"77",X"03",X"03",X"03",X"03",X"1a",X"03",X"19",X"b2",X"2e",X"3c",X"98",X"f0",X"6d",X"f0",X"6d",X"f0",X"3f",X"54",X"4d",X"d6",X"3c",X"9e",X"7c",X"5f",X"a7",X"89",X"0c",X"d6",X"d6",X"d6",X"2e",X"2e",X"1b",X"d6",X"1b",X"0b",X"3c",X"0b",X"af",X"6f",X"f3",X"f3",X"f3",X"ae",X"ae",X"82",X"d1",X"82",X"39",X"d1",X"39",X"d1",X"ff",X"d1",X"d1",X"f3",X"0b",X"3c",X"6f",X"ae",X"82",X"f3",X"22",X"f3",X"af",X"8b",X"1b",X"3c",X"0b",X"0b",X"3c",X"2e",X"98",X"2e",X"0b",X"00",X"0b",X"f3",X"ae",X"39",X"ae",X"39",X"39",X"1f",X"d1",X"d1",X"57",X"d1",X"39",X"39",X"d1",X"82",X"39",X"ae",X"0b",X"1b",X"0b",X"00",X"2e",X"2e",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"75",X"03",X"03",X"1a",X"03",X"b2",X"27",X"03",X"03",X"1a",X"00",X"00",X"f4",X"3c",X"8f",X"3c",X"8f",X"a4",X"3c",X"82",X"3c",X"a4",X"8f",X"a4",X"8f",X"a4",X"8f",X"a4",X"3c",X"82",X"3c",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",X"60",X"aa",X"aa",X"9e",X"98",X"0b",X"0b",X"1b",X"03",X"1a",X"03",X"2e",X"2f",X"62",X"62",X"15",X"cf",X"62",X"51",X"62",X"15",X"62",X"f5",X"62",X"15",X"62",X"62",X"62",X"62",X"cf",X"62",X"51",X"62",X"51",X"62",X"62",X"cf",X"15",X"62",X"62",X"62",X"62",X"62",X"51",X"77",X"62",X"51",X"62",X"51",X"62",X"51",X"cf",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"f5",X"cf",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"cf",X"62",X"ed",X"62",X"51",X"62",X"cf",X"62",X"51",X"15",X"cf",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"15",X"62",X"51",X"62",X"15",X"51",X"62",X"ed",X"2e",X"03",X"b2",X"1b",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"aa",X"84",X"0b",X"0b",X"1b",X"f0",X"03",X"1a",X"b2",X"19",X"71",X"19",X"71",X"03",X"2e",X"1b",X"6d",X"f0",X"3f",X"6d",X"f0",X"6d",X"1b",X"0b",X"ea",X"73",X"3c",X"aa",X"aa",X"a7",X"0c",X"0c",X"d6",X"d6",X"d6",X"2e",X"2e",X"2f",X"14",X"4d",X"1b",X"3c",X"8b",X"af",X"6f",X"f3",X"f3",X"f3",X"ae",X"f3",X"ae",X"ae",X"82",X"39",X"d1",X"39",X"d1",X"57",X"d1",X"39",X"d1",X"39",X"f3",X"0b",X"1b",X"0b",X"0b",X"eb",X"f3",X"f3",X"22",X"8b",X"00",X"0b",X"0b",X"3c",X"0b",X"2e",X"33",X"6d",X"2e",X"0b",X"0b",X"00",X"82",X"ae",X"39",X"4a",X"39",X"39",X"d1",X"ff",X"d1",X"d1",X"57",X"87",X"39",X"4a",X"ae",X"82",X"ad",X"3c",X"0b",X"0b",X"00",X"0b",X"2e",X"2e",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"19",X"b2",X"19",X"00",X"00",X"fb",X"00",X"a4",X"3c",X"a4",X"a4",X"00",X"82",X"3c",X"00",X"3c",X"3c",X"3c",X"a4",X"8f",X"a4",X"00",X"82",X"3c",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"9e",X"aa",X"7c",X"61",X"0b",X"1b",X"0b",X"19",X"03",X"1a",X"2e",X"2f",X"f5",X"51",X"62",X"51",X"62",X"62",X"62",X"cf",X"62",X"15",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"cf",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"61",X"62",X"62",X"62",X"15",X"62",X"62",X"15",X"62",X"cf",X"15",X"62",X"62",X"15",X"cf",X"62",X"15",X"51",X"62",X"62",X"62",X"51",X"15",X"51",X"62",X"cf",X"62",X"62",X"51",X"62",X"62",X"15",X"53",X"62",X"62",X"51",X"15",X"62",X"62",X"62",X"62",X"15",X"62",X"62",X"cf",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"cf",X"62",X"51",X"62",X"62",X"62",X"ed",X"2e",X"03",X"19",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"7c",X"9e",X"98",X"0b",X"1b",X"0b",X"2f",X"1a",X"03",X"03",X"03",X"19",X"03",X"19",X"2e",X"00",X"54",X"f0",X"6d",X"54",X"6d",X"f0",X"6d",X"f0",X"54",X"1b",X"98",X"2f",X"60",X"36",X"68",X"0c",X"89",X"d6",X"d6",X"2e",X"2e",X"d6",X"1b",X"fc",X"0b",X"0b",X"8b",X"4e",X"8b",X"af",X"4e",X"f3",X"f3",X"f3",X"ae",X"82",X"70",X"d1",X"82",X"39",X"4a",X"39",X"d1",X"57",X"d1",X"39",X"fb",X"39",X"f3",X"0b",X"3c",X"0b",X"0b",X"00",X"0b",X"eb",X"8b",X"1b",X"0b",X"0b",X"00",X"0b",X"2e",X"60",X"6d",X"93",X"2e",X"1b",X"0b",X"0b",X"39",X"ae",X"39",X"d1",X"d1",X"39",X"d1",X"d1",X"57",X"4a",X"57",X"39",X"ae",X"39",X"ae",X"82",X"ad",X"1b",X"0b",X"3c",X"0b",X"00",X"0b",X"2e",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"03",X"03",X"00",X"00",X"f4",X"3c",X"8f",X"3c",X"f4",X"8f",X"3c",X"82",X"3c",X"8f",X"a4",X"3c",X"a4",X"8f",X"a4",X"a4",X"3c",X"82",X"3c",X"f4",X"3c",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"79",X"6d",X"3f",X"6d",X"aa",X"7c",X"9e",X"aa",X"98",X"0b",X"0b",X"0b",X"03",X"b2",X"03",X"2e",X"2f",X"62",X"15",X"f5",X"62",X"15",X"f5",X"51",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"cf",X"62",X"62",X"15",X"62",X"62",X"77",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"51",X"62",X"15",X"f5",X"51",X"62",X"51",X"79",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"f5",X"62",X"62",X"15",X"62",X"15",X"cf",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"62",X"cf",X"15",X"62",X"61",X"2e",X"03",X"b2",X"1b",X"0b",X"0b",X"3b",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"79",X"03",X"03",X"b2",X"19",X"b2",X"03",X"b2",X"2e",X"1b",X"6d",X"f0",X"6d",X"3f",X"f0",X"6d",X"6d",X"aa",X"9e",X"aa",X"54",X"1b",X"aa",X"a7",X"0c",X"0c",X"a7",X"0b",X"3c",X"0b",X"0c",X"0b",X"3c",X"4d",X"1b",X"7d",X"65",X"8b",X"af",X"6f",X"f3",X"4e",X"f3",X"ae",X"f3",X"ae",X"ae",X"82",X"d1",X"39",X"d1",X"d1",X"39",X"d1",X"d1",X"57",X"39",X"d1",X"d1",X"82",X"0b",X"1b",X"0b",X"0b",X"00",X"0b",X"3c",X"0b",X"3c",X"1b",X"0b",X"2e",X"60",X"60",X"93",X"6a",X"6d",X"2e",X"0b",X"3c",X"0b",X"f3",X"4a",X"39",X"d1",X"d1",X"ff",X"d1",X"d1",X"ff",X"39",X"fb",X"39",X"ae",X"82",X"ae",X"f3",X"0b",X"0b",X"1b",X"0b",X"0b",X"3c",X"0b",X"3c",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"00",X"00",X"fb",X"00",X"a4",X"4f",X"3c",X"f4",X"3c",X"82",X"3c",X"a4",X"3c",X"a4",X"8f",X"a4",X"a4",X"8f",X"3c",X"82",X"3c",X"f4",X"3c",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",X"12",X"aa",X"aa",X"9e",X"98",X"0b",X"1b",X"0b",X"d8",X"75",X"03",X"2e",X"2f",X"62",X"62",X"51",X"62",X"cf",X"15",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"62",X"51",X"f0",X"62",X"15",X"62",X"cf",X"62",X"15",X"62",X"62",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"15",X"cf",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"62",X"62",X"62",X"79",X"62",X"62",X"62",X"15",X"cf",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"15",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"28",X"2e",X"03",X"19",X"1b",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"9e",X"98",X"0b",X"0b",X"0b",X"79",X"03",X"1a",X"03",X"03",X"03",X"19",X"03",X"e5",X"3c",X"54",X"3f",X"6d",X"f0",X"6d",X"3f",X"aa",X"7c",X"aa",X"7c",X"aa",X"60",X"a7",X"5f",X"68",X"1b",X"0b",X"ea",X"fc",X"54",X"1b",X"0b",X"2f",X"73",X"3c",X"7d",X"8b",X"4e",X"8b",X"4e",X"8b",X"f3",X"22",X"f3",X"ae",X"ae",X"70",X"d1",X"82",X"39",X"39",X"fb",X"d1",X"d1",X"57",X"d1",X"d1",X"39",X"39",X"39",X"ae",X"8b",X"1b",X"0b",X"1b",X"0b",X"0b",X"3c",X"0b",X"2e",X"2e",X"03",X"16",X"60",X"60",X"60",X"08",X"6a",X"2e",X"1b",X"0b",X"00",X"f3",X"39",X"d1",X"39",X"d1",X"57",X"d1",X"39",X"d1",X"39",X"d1",X"39",X"ae",X"ae",X"82",X"82",X"f3",X"0b",X"1b",X"0b",X"00",X"0b",X"0b",X"2e",X"2e",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"00",X"00",X"f4",X"3c",X"8f",X"4f",X"f4",X"00",X"00",X"82",X"82",X"3c",X"8f",X"a4",X"8f",X"a4",X"8f",X"3c",X"70",X"f3",X"00",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"2c",X"aa",X"7c",X"61",X"0b",X"0b",X"1b",X"19",X"71",X"03",X"2e",X"75",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"cf",X"15",X"62",X"51",X"62",X"cf",X"62",X"15",X"62",X"51",X"62",X"cf",X"15",X"f5",X"15",X"62",X"51",X"62",X"62",X"cf",X"62",X"51",X"15",X"28",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"cf",X"15",X"62",X"cf",X"62",X"62",X"15",X"51",X"62",X"62",X"51",X"62",X"cf",X"15",X"f5",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"51",X"15",X"75",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"cf",X"15",X"62",X"62",X"15",X"51",X"f5",X"cf",X"62",X"62",X"62",X"62",X"62",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"28",X"2e",X"03",X"b2",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"60",X"aa",X"98",X"0b",X"1b",X"0b",X"79",X"b2",X"03",X"19",X"71",X"19",X"b2",X"03",X"2e",X"d6",X"1b",X"0b",X"2f",X"6d",X"f0",X"6d",X"aa",X"9e",X"aa",X"9e",X"aa",X"a7",X"36",X"68",X"0c",X"0c",X"0b",X"0b",X"ea",X"fc",X"ea",X"42",X"f0",X"4d",X"e9",X"3c",X"0b",X"65",X"af",X"8b",X"f3",X"6f",X"f3",X"ae",X"f3",X"ae",X"82",X"ae",X"39",X"fb",X"39",X"57",X"39",X"d1",X"ff",X"d1",X"d1",X"d1",X"fb",X"ae",X"39",X"ae",X"82",X"8b",X"0b",X"3c",X"0b",X"3c",X"0b",X"3c",X"0b",X"2e",X"92",X"92",X"92",X"60",X"60",X"98",X"83",X"2e",X"0b",X"0b",X"0b",X"3c",X"b8",X"57",X"d1",X"d1",X"d1",X"ff",X"39",X"fb",X"39",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"f3",X"22",X"1b",X"0b",X"0b",X"00",X"0b",X"3c",X"2e",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"00",X"00",X"fb",X"00",X"a4",X"4f",X"f4",X"fb",X"f4",X"00",X"82",X"70",X"3c",X"3c",X"3c",X"3c",X"3c",X"f3",X"82",X"3c",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"12",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"cc",X"b2",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"cf",X"15",X"62",X"51",X"62",X"cf",X"62",X"62",X"51",X"62",X"62",X"15",X"cf",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"62",X"19",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"cf",X"62",X"51",X"62",X"15",X"f5",X"51",X"62",X"62",X"1a",X"15",X"62",X"15",X"f5",X"62",X"51",X"62",X"51",X"62",X"51",X"cf",X"62",X"62",X"15",X"62",X"51",X"cf",X"15",X"51",X"62",X"51",X"62",X"51",X"62",X"cf",X"15",X"62",X"51",X"62",X"62",X"15",X"75",X"2e",X"19",X"03",X"0b",X"0b",X"1b",X"17",X"3f",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"33",X"0b",X"0b",X"1b",X"2f",X"03",X"19",X"71",X"19",X"03",X"03",X"2e",X"1b",X"0b",X"2e",X"4d",X"1b",X"0b",X"54",X"f0",X"60",X"aa",X"7c",X"aa",X"6d",X"a7",X"a7",X"0c",X"0c",X"d6",X"d6",X"0c",X"1b",X"0b",X"ea",X"42",X"f0",X"14",X"e9",X"3c",X"1b",X"8b",X"4e",X"8b",X"4e",X"f3",X"f3",X"f3",X"ae",X"ae",X"ae",X"39",X"ae",X"39",X"39",X"4a",X"d1",X"57",X"d1",X"57",X"d1",X"39",X"39",X"39",X"ae",X"ae",X"f3",X"ae",X"82",X"6f",X"1b",X"0b",X"0b",X"0b",X"3c",X"0b",X"2e",X"69",X"92",X"69",X"92",X"33",X"60",X"60",X"2e",X"1b",X"3c",X"0b",X"0b",X"f3",X"d1",X"ff",X"d1",X"39",X"1f",X"39",X"39",X"39",X"ae",X"82",X"ae",X"f3",X"f3",X"22",X"48",X"f3",X"4e",X"1b",X"0b",X"0b",X"3c",X"0b",X"ec",X"27",X"19",X"b2",X"03",X"03",X"19",X"b2",X"19",X"03",X"19",X"03",X"1a",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"fb",X"f4",X"91",X"00",X"00",X"82",X"82",X"70",X"82",X"82",X"82",X"70",X"3c",X"00",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"cd",X"6d",X"f0",X"6d",X"f0",X"60",X"aa",X"aa",X"92",X"61",X"0b",X"0b",X"0b",X"19",X"03",X"75",X"03",X"2e",X"1a",X"15",X"f5",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"15",X"75",X"2e",X"1a",X"15",X"f5",X"51",X"62",X"62",X"51",X"15",X"62",X"62",X"15",X"62",X"62",X"15",X"62",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"62",X"51",X"62",X"62",X"28",X"2e",X"1a",X"62",X"51",X"62",X"15",X"51",X"62",X"62",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"62",X"62",X"15",X"62",X"62",X"15",X"62",X"51",X"62",X"15",X"f5",X"51",X"1a",X"2e",X"03",X"b2",X"03",X"0b",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"9e",X"aa",X"7c",X"61",X"0b",X"0b",X"0b",X"79",X"03",X"b2",X"19",X"03",X"1a",X"ec",X"0b",X"0b",X"2f",X"0b",X"1b",X"42",X"fc",X"2f",X"0b",X"3c",X"aa",X"aa",X"9e",X"a7",X"5f",X"89",X"0c",X"f8",X"d6",X"2e",X"2e",X"d6",X"1b",X"3c",X"f0",X"fc",X"54",X"4d",X"e9",X"00",X"0b",X"65",X"8b",X"f3",X"4e",X"f3",X"ae",X"f3",X"ae",X"70",X"ae",X"39",X"39",X"fb",X"57",X"39",X"d1",X"d1",X"d1",X"39",X"1f",X"39",X"ae",X"39",X"ae",X"82",X"f3",X"22",X"f3",X"f3",X"4e",X"8b",X"3c",X"0b",X"0b",X"3c",X"2e",X"c3",X"2e",X"2e",X"ec",X"69",X"60",X"60",X"2e",X"2e",X"3c",X"0b",X"3c",X"38",X"f3",X"ff",X"d1",X"39",X"39",X"4a",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"f3",X"f3",X"6f",X"8b",X"3c",X"0b",X"3c",X"0b",X"0b",X"2e",X"03",X"b2",X"03",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"00",X"00",X"fb",X"00",X"a4",X"4f",X"f4",X"fb",X"f4",X"fb",X"f4",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"fb",X"f4",X"fb",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"aa",X"60",X"aa",X"98",X"0b",X"0b",X"7d",X"03",X"b2",X"27",X"03",X"30",X"19",X"1a",X"15",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"51",X"62",X"15",X"f5",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"15",X"62",X"51",X"62",X"62",X"51",X"19",X"b2",X"2e",X"03",X"1a",X"15",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"51",X"62",X"51",X"15",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"1a",X"03",X"cc",X"03",X"1a",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"15",X"1a",X"03",X"cc",X"03",X"03",X"19",X"0b",X"0b",X"0b",X"61",X"f0",X"6d",X"6d",X"f0",
    X"aa",X"7c",X"0d",X"9e",X"98",X"0b",X"1b",X"83",X"2f",X"19",X"03",X"03",X"b2",X"03",X"2e",X"0b",X"2f",X"6d",X"f0",X"54",X"3c",X"0b",X"ea",X"42",X"fc",X"54",X"e4",X"54",X"36",X"a7",X"0c",X"0c",X"d6",X"d6",X"2e",X"2e",X"0c",X"0b",X"d6",X"6d",X"4d",X"3f",X"ea",X"e9",X"3c",X"1b",X"0b",X"af",X"65",X"f3",X"f3",X"f3",X"ae",X"82",X"ae",X"39",X"ae",X"39",X"39",X"fb",X"57",X"d1",X"57",X"d1",X"57",X"39",X"d1",X"39",X"ae",X"82",X"82",X"ae",X"f3",X"f3",X"8b",X"4e",X"8b",X"3c",X"0b",X"3c",X"0b",X"30",X"2e",X"1b",X"0b",X"0b",X"2e",X"ec",X"2e",X"60",X"60",X"2e",X"1b",X"0b",X"0b",X"3c",X"b8",X"39",X"1f",X"39",X"d1",X"39",X"ae",X"ae",X"82",X"82",X"f3",X"f3",X"4e",X"f3",X"af",X"0b",X"0b",X"0b",X"3c",X"3c",X"2e",X"19",X"03",X"75",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"91",X"f4",X"fb",X"f4",X"91",X"f4",X"fb",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"92",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"d8",X"1a",X"03",X"b2",X"03",X"2e",X"03",X"75",X"75",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"51",X"75",X"03",X"1a",X"ec",X"03",X"2e",X"19",X"1a",X"75",X"15",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"15",X"51",X"75",X"75",X"03",X"cc",X"03",X"21",X"03",X"1a",X"75",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"15",X"51",X"75",X"75",X"03",X"2e",X"03",X"1a",X"03",X"b2",X"1b",X"0b",X"0b",X"3b",X"6d",X"f0",X"3f",X"6d",
    X"9e",X"aa",X"7c",X"aa",X"98",X"1b",X"0b",X"1b",X"2f",X"03",X"b2",X"03",X"1a",X"03",X"2e",X"0b",X"f0",X"6d",X"3f",X"6d",X"f0",X"54",X"1b",X"f0",X"ea",X"42",X"ea",X"f0",X"0b",X"3c",X"68",X"0c",X"d6",X"2e",X"2e",X"2e",X"aa",X"1b",X"d6",X"fc",X"54",X"fc",X"54",X"4d",X"e9",X"ab",X"0b",X"0b",X"f3",X"6f",X"f3",X"ae",X"f3",X"ae",X"ae",X"ae",X"39",X"fb",X"39",X"d1",X"39",X"d1",X"d1",X"57",X"b8",X"d1",X"39",X"ae",X"39",X"ae",X"82",X"f3",X"f3",X"4e",X"f3",X"4e",X"8b",X"0b",X"3c",X"0b",X"0b",X"0b",X"0b",X"3c",X"0b",X"1b",X"0b",X"0b",X"0b",X"2e",X"2e",X"ec",X"2e",X"3c",X"0b",X"0b",X"3c",X"8b",X"39",X"39",X"4a",X"82",X"39",X"ae",X"f3",X"ae",X"f3",X"22",X"f3",X"6f",X"8b",X"4e",X"0b",X"00",X"0b",X"0b",X"2e",X"03",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"00",X"00",X"fb",X"00",X"a4",X"91",X"f4",X"fb",X"f4",X"91",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"79",X"6d",X"f0",X"60",X"aa",X"aa",X"60",X"61",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"03",X"03",X"b2",X"2e",X"2e",X"03",X"1a",X"75",X"1a",X"f0",X"f0",X"98",X"f0",X"f0",X"98",X"f0",X"f0",X"ed",X"f0",X"54",X"f0",X"2f",X"f0",X"f0",X"54",X"28",X"f0",X"1a",X"19",X"03",X"1a",X"2e",X"03",X"19",X"71",X"30",X"2e",X"19",X"19",X"75",X"28",X"f0",X"f0",X"61",X"79",X"61",X"79",X"79",X"61",X"79",X"61",X"77",X"2f",X"f0",X"2f",X"f0",X"61",X"f0",X"79",X"1a",X"19",X"03",X"21",X"2e",X"03",X"1a",X"03",X"21",X"03",X"03",X"1a",X"1a",X"28",X"f0",X"f0",X"98",X"2f",X"f0",X"98",X"f0",X"f0",X"f0",X"ed",X"f0",X"f0",X"f0",X"98",X"f0",X"f0",X"f0",X"f0",X"1a",X"19",X"03",X"2e",X"2e",X"1a",X"03",X"b2",X"03",X"19",X"3c",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"9e",X"54",X"0b",X"0b",X"0b",X"ed",X"03",X"19",X"1a",X"03",X"2e",X"3c",X"54",X"f0",X"6d",X"f0",X"6d",X"f0",X"0b",X"d6",X"d6",X"98",X"f0",X"42",X"ea",X"42",X"f0",X"3c",X"0b",X"d6",X"2e",X"2e",X"d6",X"1b",X"73",X"32",X"32",X"3f",X"4d",X"aa",X"42",X"e9",X"4d",X"1b",X"3c",X"0b",X"f3",X"f3",X"f3",X"ae",X"ae",X"70",X"39",X"ae",X"39",X"39",X"d1",X"d1",X"d1",X"ff",X"d1",X"0b",X"1b",X"0b",X"b8",X"ae",X"ae",X"f3",X"ae",X"f3",X"f3",X"6f",X"8b",X"af",X"0b",X"00",X"0b",X"3c",X"0b",X"3c",X"1b",X"0b",X"3c",X"0b",X"1b",X"0b",X"3c",X"0b",X"0b",X"0b",X"3c",X"2e",X"3c",X"0b",X"3c",X"0b",X"4e",X"39",X"d1",X"82",X"ae",X"ae",X"f3",X"f3",X"f3",X"48",X"f3",X"4e",X"8b",X"1b",X"0b",X"0b",X"00",X"0b",X"2e",X"03",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"71",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f4",X"fb",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"f4",X"fb",X"f4",X"fb",X"f4",X"91",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"aa",X"92",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"2e",X"2e",X"2e",X"ec",X"2e",X"2e",X"ec",X"2e",X"2e",X"ec",X"2e",X"2e",X"2e",X"2e",X"ec",X"2e",X"2e",X"2e",X"2e",X"30",X"2e",X"2e",X"ec",X"2e",X"2e",X"2e",X"03",X"b2",X"03",X"e5",X"03",X"75",X"75",X"51",X"62",X"62",X"cf",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"cf",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"19",X"75",X"03",X"2e",X"03",X"03",X"1a",X"2e",X"2e",X"ec",X"2e",X"2e",X"2e",X"ec",X"2e",X"e5",X"2e",X"ec",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"2e",X"2e",X"ec",X"2e",X"2e",X"2e",X"2e",X"b2",X"19",X"03",X"03",X"19",X"03",X"b2",X"ad",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"84",X"0b",X"1b",X"0b",X"79",X"03",X"b2",X"03",X"03",X"e5",X"0b",X"f0",X"6d",X"f0",X"6d",X"3f",X"54",X"f0",X"4d",X"d6",X"d6",X"fc",X"2f",X"42",X"fc",X"42",X"ea",X"54",X"1b",X"0b",X"d6",X"aa",X"0b",X"4d",X"e9",X"32",X"f0",X"4d",X"fc",X"2f",X"4d",X"e9",X"7a",X"0b",X"1b",X"0b",X"f3",X"ae",X"f3",X"82",X"ae",X"ae",X"39",X"39",X"fb",X"d1",X"39",X"d1",X"57",X"d1",X"f3",X"0b",X"3c",X"0b",X"1b",X"38",X"ae",X"f3",X"f3",X"6f",X"f3",X"af",X"6f",X"1b",X"0b",X"0b",X"0b",X"3c",X"8b",X"8b",X"f3",X"4e",X"0b",X"1b",X"0b",X"1b",X"3c",X"0b",X"3c",X"0b",X"1b",X"0b",X"0b",X"0b",X"3c",X"0b",X"3c",X"eb",X"39",X"ae",X"82",X"ae",X"f3",X"f3",X"22",X"af",X"8b",X"af",X"0b",X"1b",X"0b",X"0b",X"3c",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"19",X"03",X"1a",X"03",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"4f",X"fb",X"91",X"f4",X"4f",X"fb",X"f4",X"fb",X"f4",X"4f",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"60",X"aa",X"aa",X"84",X"0b",X"0b",X"0b",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"19",X"71",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"b2",X"03",X"03",X"19",X"21",X"03",X"75",X"62",X"62",X"62",X"51",X"62",X"51",X"f5",X"62",X"62",X"15",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"51",X"cf",X"15",X"62",X"51",X"62",X"75",X"19",X"ec",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"b2",X"27",X"19",X"1b",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"3f",
    X"9e",X"aa",X"60",X"aa",X"98",X"0b",X"0b",X"1b",X"2f",X"03",X"1a",X"03",X"cc",X"0b",X"2f",X"6d",X"3f",X"6d",X"f0",X"6d",X"1b",X"f0",X"73",X"3c",X"1b",X"54",X"ea",X"54",X"f0",X"ea",X"fc",X"ea",X"fc",X"2f",X"0b",X"0b",X"42",X"bc",X"14",X"e9",X"32",X"3f",X"14",X"2f",X"73",X"e9",X"00",X"ae",X"0b",X"3c",X"0b",X"f3",X"ae",X"ae",X"ae",X"39",X"ae",X"39",X"39",X"39",X"1f",X"57",X"d1",X"d1",X"ff",X"f3",X"0b",X"1b",X"0b",X"3c",X"0b",X"3c",X"eb",X"f3",X"22",X"8b",X"af",X"0b",X"1b",X"0b",X"3c",X"0b",X"eb",X"4e",X"8b",X"f3",X"22",X"70",X"6f",X"0b",X"0b",X"0b",X"1b",X"0b",X"00",X"0b",X"0b",X"00",X"0b",X"0b",X"0b",X"0b",X"00",X"65",X"ae",X"f3",X"ae",X"f3",X"f3",X"f3",X"8b",X"4e",X"0b",X"3c",X"0b",X"3c",X"0b",X"2e",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"19",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f4",X"f4",X"f4",X"f4",X"fb",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"f4",X"fb",X"f4",X"fb",X"f4",X"3c",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"9e",X"aa",X"aa",X"7c",X"61",X"0b",X"0b",X"1b",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"b2",X"2e",X"03",X"28",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"15",X"51",X"cf",X"62",X"62",X"62",X"51",X"62",X"cf",X"62",X"15",X"51",X"62",X"cf",X"15",X"62",X"62",X"62",X"cf",X"15",X"62",X"62",X"28",X"2e",X"03",X"03",X"19",X"03",X"b2",X"27",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"b2",X"83",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"9e",X"98",X"0b",X"1b",X"83",X"2f",X"03",X"03",X"03",X"e5",X"1b",X"6d",X"f0",X"6d",X"f0",X"6d",X"2f",X"98",X"ea",X"73",X"2f",X"9e",X"7c",X"2f",X"0b",X"d6",X"54",X"1b",X"0b",X"0b",X"ea",X"42",X"fc",X"2f",X"42",X"ea",X"73",X"4d",X"1b",X"0b",X"1b",X"ea",X"14",X"1b",X"82",X"ae",X"0b",X"0b",X"1b",X"82",X"ae",X"70",X"ae",X"d1",X"39",X"fb",X"57",X"39",X"d1",X"d1",X"57",X"39",X"1f",X"22",X"8b",X"3c",X"0b",X"0b",X"0b",X"00",X"0b",X"3c",X"8b",X"4e",X"0b",X"2e",X"3c",X"0b",X"0b",X"af",X"8b",X"f3",X"6f",X"f3",X"22",X"ae",X"70",X"39",X"ae",X"f3",X"0b",X"0b",X"1b",X"3c",X"0b",X"0b",X"00",X"0b",X"1b",X"0b",X"0b",X"af",X"ae",X"f3",X"22",X"f3",X"4e",X"f3",X"6f",X"3c",X"0b",X"0b",X"3c",X"0b",X"ec",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"19",X"03",X"1a",X"03",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"fb",X"82",X"70",X"f3",X"82",X"70",X"82",X"82",X"70",X"82",X"82",X"70",X"f3",X"f4",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"6d",X"aa",X"7c",X"0d",X"9e",X"98",X"0b",X"1b",X"0b",X"d8",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"75",X"03",X"b2",X"03",X"2e",X"19",X"15",X"f5",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"62",X"cf",X"15",X"62",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"19",X"21",X"03",X"b2",X"d8",X"19",X"71",X"75",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"71",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"19",X"03",X"19",X"03",X"1a",X"03",X"b2",X"19",X"3c",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"9e",X"aa",X"7c",X"61",X"0b",X"0b",X"1b",X"2f",X"19",X"b2",X"2e",X"3c",X"0b",X"f0",X"6d",X"3f",X"6d",X"f0",X"0b",X"6d",X"fc",X"6d",X"2f",X"a7",X"36",X"9e",X"1b",X"d6",X"d6",X"54",X"0c",X"a7",X"0b",X"3c",X"0b",X"d6",X"98",X"fc",X"ea",X"4d",X"1b",X"82",X"48",X"0b",X"0b",X"1b",X"82",X"b7",X"82",X"ad",X"3c",X"0b",X"82",X"ae",X"39",X"ae",X"39",X"39",X"4a",X"d1",X"57",X"ff",X"d1",X"d1",X"39",X"39",X"39",X"6f",X"1b",X"0b",X"3c",X"0b",X"0b",X"0b",X"3c",X"0b",X"ec",X"2e",X"1b",X"0b",X"00",X"8b",X"4e",X"af",X"f3",X"f3",X"ae",X"f3",X"ae",X"ae",X"39",X"d1",X"39",X"39",X"22",X"0b",X"0b",X"1b",X"0b",X"0b",X"3c",X"1b",X"0b",X"0b",X"00",X"8b",X"f3",X"f3",X"22",X"8b",X"af",X"0b",X"0b",X"3c",X"0b",X"0b",X"2e",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"70",X"f4",X"91",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"53",X"79",X"6d",X"0d",X"f0",X"9e",X"aa",X"7c",X"aa",X"23",X"0b",X"0b",X"0b",X"19",X"03",X"75",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"27",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"71",X"03",X"03",X"b2",X"03",X"19",X"03",X"cc",X"1a",X"51",X"62",X"62",X"cf",X"15",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"f5",X"62",X"51",X"15",X"62",X"62",X"28",X"2e",X"03",X"19",X"b2",X"27",X"19",X"03",X"03",X"b2",X"19",X"71",X"19",X"03",X"03",X"b2",X"27",X"19",X"03",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"0b",X"0b",X"0b",X"17",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"0d",X"aa",X"33",X"0b",X"0b",X"0b",X"ed",X"03",X"03",X"2e",X"0b",X"ed",X"6d",X"f0",X"6d",X"f0",X"54",X"0b",X"2f",X"42",X"2f",X"6d",X"5f",X"a7",X"54",X"f0",X"e9",X"2f",X"aa",X"d6",X"2e",X"d6",X"a7",X"3c",X"d6",X"d6",X"f0",X"42",X"fc",X"0b",X"ae",X"82",X"ae",X"ae",X"8b",X"ae",X"82",X"ae",X"82",X"0b",X"1b",X"0b",X"65",X"82",X"39",X"39",X"4a",X"57",X"39",X"d1",X"d1",X"d1",X"39",X"ff",X"39",X"fb",X"ae",X"39",X"8b",X"1b",X"1b",X"0b",X"00",X"0b",X"0b",X"2e",X"2e",X"3c",X"0b",X"0b",X"eb",X"8b",X"f3",X"4e",X"f3",X"f3",X"ae",X"ae",X"39",X"ae",X"39",X"39",X"4a",X"39",X"d1",X"57",X"d1",X"ae",X"f3",X"0b",X"0b",X"0b",X"1b",X"0b",X"00",X"0b",X"0b",X"65",X"f3",X"6f",X"3c",X"0b",X"3c",X"0b",X"30",X"03",X"1a",X"03",X"03",X"19",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"6d",X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"2e",X"28",X"62",X"15",X"51",X"62",X"62",X"cf",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"15",X"cf",X"15",X"f5",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"cf",X"62",X"2f",X"2e",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"1a",X"71",X"75",X"03",X"03",X"b2",X"03",X"19",X"b2",X"27",X"19",X"03",X"1a",X"03",X"19",X"71",X"03",X"19",X"03",X"75",X"03",X"03",X"b2",X"19",X"1b",X"0b",X"3c",X"33",X"f0",X"6d",X"3f",X"6d",
    X"9e",X"aa",X"7c",X"aa",X"98",X"0b",X"1b",X"0b",X"79",X"03",X"1a",X"2e",X"3c",X"6d",X"f0",X"6d",X"f0",X"6d",X"9e",X"aa",X"7c",X"f0",X"0b",X"5f",X"a7",X"6d",X"1b",X"42",X"bc",X"1b",X"d6",X"2e",X"2e",X"a7",X"3c",X"73",X"4d",X"1b",X"0b",X"1b",X"0b",X"0b",X"82",X"ae",X"70",X"ae",X"82",X"ae",X"82",X"b7",X"82",X"ae",X"48",X"0b",X"1b",X"0b",X"ae",X"39",X"d1",X"87",X"d1",X"57",X"d1",X"57",X"d1",X"39",X"4a",X"39",X"39",X"ae",X"ae",X"f3",X"8b",X"1b",X"0b",X"00",X"0b",X"00",X"0b",X"3c",X"0b",X"3c",X"8b",X"4e",X"8b",X"f3",X"f3",X"ae",X"f3",X"ae",X"ae",X"39",X"39",X"fb",X"39",X"d1",X"d1",X"d1",X"d1",X"39",X"d1",X"39",X"ae",X"39",X"ae",X"48",X"0b",X"0b",X"1b",X"0b",X"0b",X"00",X"0b",X"0b",X"0b",X"3c",X"0b",X"2e",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"33",X"f0",X"6d",X"6d",X"f0",X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"19",X"03",X"19",X"03",X"75",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"cc",X"54",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"cf",X"15",X"62",X"15",X"62",X"51",X"62",X"cf",X"15",X"62",X"51",X"62",X"62",X"62",X"15",X"62",X"cf",X"62",X"15",X"62",X"62",X"51",X"15",X"f5",X"2f",X"2e",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"75",X"03",X"b2",X"19",X"03",X"03",X"19",X"b2",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"0b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"60",X"61",X"0b",X"0b",X"0b",X"2f",X"03",X"e5",X"1b",X"0b",X"f0",X"6d",X"3f",X"6d",X"f0",X"aa",X"2c",X"aa",X"aa",X"6d",X"36",X"a7",X"0b",X"2f",X"42",X"fc",X"0b",X"d6",X"2e",X"2e",X"aa",X"0b",X"4d",X"e9",X"3c",X"ae",X"8b",X"0b",X"7d",X"ae",X"82",X"ae",X"82",X"b7",X"82",X"ae",X"82",X"ae",X"82",X"ae",X"82",X"ad",X"3c",X"0b",X"eb",X"39",X"ff",X"39",X"d1",X"57",X"d1",X"d1",X"d1",X"39",X"d1",X"82",X"39",X"ae",X"ae",X"f3",X"f3",X"6f",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"3c",X"6f",X"af",X"f3",X"6f",X"f3",X"f3",X"ae",X"82",X"39",X"ae",X"39",X"39",X"d1",X"39",X"d1",X"d1",X"57",X"d1",X"39",X"d1",X"39",X"ae",X"82",X"f3",X"ae",X"f3",X"82",X"8b",X"1b",X"0b",X"3c",X"0b",X"00",X"0b",X"0b",X"3c",X"2e",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"71",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"70",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"3b",X"6d",X"f0",X"3f",X"f0",X"60",X"aa",X"aa",X"9e",X"98",X"0b",X"0b",X"7d",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"27",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"2e",X"ed",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"cf",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"03",X"19",X"03",X"19",X"71",X"19",X"3c",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"28",X"03",X"2e",X"00",X"0b",X"2f",X"6d",X"f0",X"6d",X"aa",X"12",X"aa",X"9e",X"aa",X"7c",X"5f",X"a7",X"aa",X"0b",X"0b",X"3c",X"d6",X"2e",X"2e",X"d6",X"1b",X"42",X"ea",X"14",X"1b",X"ae",X"70",X"ae",X"48",X"82",X"b7",X"82",X"ae",X"82",X"ae",X"ae",X"82",X"ae",X"ae",X"ae",X"82",X"ae",X"8b",X"0b",X"00",X"8b",X"eb",X"d1",X"d1",X"d1",X"d1",X"d1",X"39",X"39",X"4a",X"39",X"ae",X"82",X"f3",X"ae",X"f3",X"82",X"4e",X"4e",X"0b",X"3c",X"0b",X"3c",X"0b",X"eb",X"8b",X"4e",X"f3",X"f3",X"82",X"f3",X"ae",X"ae",X"39",X"d1",X"4a",X"39",X"d1",X"39",X"ff",X"d1",X"d1",X"d1",X"39",X"ae",X"39",X"ae",X"ae",X"f3",X"f3",X"22",X"4e",X"f3",X"8b",X"4e",X"1b",X"0b",X"0b",X"3c",X"0b",X"2e",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"6d",X"aa",X"12",X"aa",X"7c",X"61",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"19",X"71",X"19",X"71",X"19",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"2e",X"2f",X"62",X"51",X"62",X"15",X"f5",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"15",X"62",X"cf",X"15",X"62",X"62",X"62",X"51",X"79",X"2e",X"03",X"75",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"71",X"19",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"b2",X"03",X"19",X"1b",X"0b",X"1b",X"3b",X"6d",X"f0",X"3f",X"6d",
    X"9e",X"aa",X"aa",X"12",X"98",X"1b",X"0b",X"0b",X"79",X"1a",X"2e",X"2e",X"1b",X"0b",X"00",X"54",X"f0",X"9e",X"aa",X"7c",X"aa",X"6d",X"9e",X"a7",X"0c",X"68",X"0c",X"aa",X"0b",X"d6",X"2e",X"ec",X"a7",X"0b",X"ea",X"fc",X"42",X"0b",X"ae",X"82",X"ae",X"82",X"ae",X"82",X"ae",X"82",X"ae",X"39",X"39",X"d1",X"39",X"39",X"4a",X"39",X"57",X"39",X"ae",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"0b",X"1b",X"0b",X"0b",X"00",X"8b",X"ae",X"82",X"f3",X"22",X"8b",X"f3",X"8b",X"00",X"0b",X"0b",X"3c",X"0b",X"3c",X"8b",X"4e",X"8b",X"46",X"f3",X"ae",X"82",X"ae",X"82",X"39",X"39",X"39",X"d1",X"d1",X"d1",X"d1",X"d1",X"39",X"4a",X"39",X"ae",X"ae",X"f3",X"ae",X"f3",X"f3",X"f3",X"6f",X"af",X"8b",X"0b",X"00",X"0b",X"3c",X"0b",X"2e",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"f0",X"6d",X"6d",X"f0",X"aa",X"6d",X"aa",X"aa",X"84",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"75",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"2e",X"2f",X"62",X"62",X"cf",X"62",X"15",X"62",X"15",X"cf",X"15",X"62",X"62",X"15",X"62",X"62",X"62",X"cf",X"62",X"15",X"51",X"62",X"62",X"cf",X"62",X"51",X"62",X"51",X"62",X"cf",X"15",X"51",X"62",X"61",X"2e",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"83",X"0b",X"0b",X"98",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"9e",X"2c",X"ba",X"0b",X"1b",X"0b",X"77",X"03",X"03",X"b2",X"2e",X"2e",X"0b",X"1b",X"0b",X"00",X"54",X"aa",X"9e",X"aa",X"a7",X"36",X"68",X"0c",X"0c",X"09",X"d6",X"d6",X"2e",X"2e",X"aa",X"0b",X"fc",X"ea",X"ea",X"e4",X"82",X"ae",X"70",X"ae",X"ae",X"ae",X"39",X"d1",X"39",X"4a",X"39",X"4a",X"39",X"d1",X"57",X"d1",X"ae",X"0b",X"0b",X"3c",X"1b",X"54",X"f0",X"54",X"2f",X"54",X"2f",X"54",X"54",X"f0",X"0b",X"0b",X"1b",X"0b",X"65",X"f3",X"f3",X"6f",X"af",X"8b",X"1b",X"0b",X"00",X"0b",X"0b",X"af",X"6f",X"f3",X"8b",X"f3",X"82",X"ae",X"70",X"d1",X"82",X"d1",X"87",X"d1",X"39",X"d1",X"57",X"d1",X"ff",X"39",X"fb",X"39",X"ae",X"82",X"f3",X"f3",X"46",X"8b",X"f3",X"4e",X"8b",X"1b",X"0b",X"0b",X"0b",X"3c",X"2e",X"1a",X"03",X"19",X"71",X"03",X"1a",X"03",X"1a",X"03",X"03",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"53",X"6d",X"f0",X"3f",X"f0",X"12",X"aa",X"7c",X"9e",X"98",X"0b",X"1b",X"0b",X"03",X"b2",X"27",X"1a",X"03",X"71",X"27",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"19",X"03",X"71",X"2e",X"ed",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"cf",X"15",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"15",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"15",X"61",X"2e",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"75",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"b2",X"27",X"19",X"3c",X"0b",X"1b",X"3b",X"f0",X"6d",X"3f",X"6d",
    X"9e",X"aa",X"aa",X"aa",X"98",X"0b",X"0b",X"0b",X"2f",X"03",X"06",X"19",X"03",X"03",X"cc",X"2e",X"3c",X"0b",X"0b",X"1b",X"0b",X"2f",X"a7",X"68",X"0c",X"0c",X"f8",X"d6",X"d6",X"2e",X"2e",X"2e",X"3c",X"0b",X"0b",X"0b",X"0b",X"0b",X"82",X"ae",X"ae",X"ae",X"39",X"4a",X"39",X"4a",X"39",X"d1",X"39",X"39",X"d1",X"57",X"ae",X"0b",X"3c",X"54",X"f0",X"54",X"54",X"2f",X"54",X"2f",X"54",X"2f",X"54",X"2f",X"54",X"2f",X"54",X"2f",X"54",X"f0",X"0b",X"3c",X"6f",X"f3",X"4e",X"8b",X"00",X"0b",X"0b",X"0b",X"00",X"eb",X"8b",X"4e",X"f3",X"22",X"ae",X"f3",X"ae",X"ae",X"39",X"39",X"39",X"d1",X"d1",X"ff",X"d1",X"d1",X"39",X"d1",X"39",X"ae",X"39",X"ae",X"ae",X"f3",X"f3",X"f3",X"4e",X"8b",X"4e",X"0b",X"3c",X"0b",X"3c",X"0b",X"2e",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"b2",X"19",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"4f",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"6d",X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"03",X"19",X"03",X"b2",X"19",X"2e",X"2f",X"62",X"15",X"62",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"62",X"15",X"62",X"62",X"51",X"cf",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"ed",X"2e",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"03",X"75",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"aa",X"92",X"aa",X"98",X"1b",X"0b",X"1b",X"61",X"03",X"03",X"03",X"e5",X"2e",X"3c",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"aa",X"0c",X"68",X"d6",X"d6",X"d6",X"2e",X"2e",X"d6",X"1b",X"0b",X"82",X"ae",X"82",X"b7",X"82",X"b7",X"82",X"39",X"d1",X"39",X"39",X"d1",X"39",X"39",X"d1",X"d1",X"ae",X"0b",X"0b",X"54",X"f0",X"54",X"2f",X"54",X"2f",X"54",X"1b",X"0b",X"0b",X"00",X"0b",X"0b",X"2f",X"54",X"2f",X"54",X"2f",X"54",X"f0",X"6d",X"3c",X"3c",X"6f",X"af",X"0b",X"0b",X"3c",X"1b",X"0b",X"0b",X"af",X"f3",X"8b",X"f3",X"f3",X"ae",X"82",X"39",X"ae",X"39",X"d1",X"d1",X"39",X"d1",X"d1",X"57",X"d1",X"d1",X"39",X"39",X"ae",X"ae",X"f3",X"ae",X"f3",X"f3",X"22",X"8b",X"af",X"8b",X"1b",X"0b",X"0b",X"00",X"0b",X"2e",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"f4",X"f4",X"3c",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"6d",X"f0",X"aa",X"7c",X"aa",X"9e",X"98",X"1b",X"0b",X"0b",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"75",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"27",X"19",X"03",X"cc",X"54",X"62",X"62",X"51",X"62",X"cf",X"15",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"f5",X"62",X"62",X"15",X"f5",X"51",X"62",X"ed",X"2e",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"71",X"19",X"03",X"1a",X"03",X"1a",X"03",X"71",X"19",X"71",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"b2",X"27",X"19",X"03",X"1a",X"03",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"60",X"aa",X"9e",X"98",X"0b",X"0b",X"0b",X"2f",X"03",X"1a",X"2e",X"2f",X"0b",X"6d",X"aa",X"9e",X"aa",X"7c",X"f0",X"0b",X"0b",X"42",X"1b",X"0b",X"aa",X"5f",X"f8",X"f8",X"2e",X"2e",X"aa",X"42",X"3c",X"f3",X"ae",X"ae",X"82",X"ae",X"82",X"ae",X"39",X"39",X"d1",X"d1",X"d1",X"d1",X"d1",X"d1",X"d1",X"0b",X"2f",X"54",X"2f",X"54",X"2f",X"54",X"2f",X"0b",X"3c",X"0b",X"3c",X"0b",X"3c",X"0b",X"3c",X"0b",X"1b",X"0b",X"00",X"54",X"ed",X"54",X"2f",X"54",X"6d",X"1b",X"8b",X"0b",X"00",X"0b",X"0b",X"0b",X"00",X"0b",X"eb",X"f3",X"22",X"ae",X"f3",X"ae",X"ae",X"39",X"39",X"4a",X"39",X"d1",X"ff",X"d1",X"d1",X"39",X"d1",X"39",X"ae",X"39",X"ae",X"82",X"f3",X"f3",X"f3",X"6f",X"f3",X"4e",X"eb",X"0b",X"1b",X"0b",X"3c",X"0b",X"2e",X"03",X"03",X"b2",X"03",X"19",X"1a",X"03",X"b2",X"19",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"f0",X"3f",X"f0",X"60",X"aa",X"aa",X"7c",X"61",X"0b",X"0b",X"1b",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"19",X"71",X"03",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"2e",X"ed",X"62",X"51",X"62",X"15",X"51",X"62",X"62",X"cf",X"62",X"15",X"62",X"15",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"54",X"2e",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"b2",X"27",X"19",X"0b",X"1b",X"0b",X"53",X"6d",X"f0",X"6d",X"3f",
    X"9e",X"aa",X"aa",X"7c",X"61",X"0b",X"1b",X"0b",X"79",X"03",X"2e",X"2f",X"0b",X"3f",X"aa",X"7c",X"aa",X"aa",X"60",X"aa",X"a7",X"2f",X"0b",X"d6",X"42",X"42",X"0b",X"1b",X"9e",X"a7",X"f8",X"0b",X"42",X"bc",X"0b",X"f3",X"82",X"ae",X"82",X"ae",X"d1",X"39",X"d1",X"d1",X"57",X"8b",X"0b",X"1b",X"0b",X"0b",X"2f",X"54",X"2f",X"54",X"2f",X"54",X"0b",X"3c",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"2f",X"54",X"2f",X"54",X"f0",X"0b",X"1b",X"0b",X"3c",X"0b",X"1b",X"0b",X"0b",X"00",X"eb",X"f3",X"f3",X"ae",X"ae",X"39",X"ae",X"d1",X"39",X"d1",X"39",X"d1",X"57",X"d1",X"ae",X"ae",X"39",X"4a",X"ae",X"82",X"82",X"ae",X"f3",X"22",X"82",X"8b",X"8b",X"4e",X"0b",X"3c",X"0b",X"0b",X"3c",X"2e",X"03",X"1a",X"03",X"19",X"71",X"03",X"03",X"19",X"03",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"f4",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"6d",X"aa",X"aa",X"60",X"aa",X"84",X"0b",X"0b",X"1b",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"ec",X"f0",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"cf",X"62",X"62",X"15",X"cf",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"cf",X"15",X"62",X"62",X"62",X"cf",X"62",X"2f",X"2e",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"0b",X"0b",X"0b",X"3b",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"9e",X"98",X"0b",X"0b",X"0b",X"79",X"2e",X"0b",X"54",X"f0",X"6d",X"aa",X"9e",X"aa",X"9e",X"aa",X"aa",X"90",X"0c",X"54",X"2f",X"d6",X"d6",X"d6",X"32",X"42",X"3c",X"3f",X"1b",X"ea",X"ea",X"42",X"1b",X"ae",X"57",X"d1",X"d1",X"39",X"d1",X"ff",X"4e",X"0b",X"2f",X"2f",X"54",X"3c",X"54",X"f0",X"54",X"2f",X"0b",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"3c",X"54",X"ed",X"54",X"6d",X"3c",X"0b",X"17",X"e4",X"0b",X"1b",X"0b",X"0b",X"f3",X"ae",X"f3",X"ae",X"82",X"39",X"39",X"39",X"4a",X"57",X"d1",X"d1",X"57",X"39",X"0b",X"3c",X"0b",X"65",X"ae",X"82",X"f3",X"f3",X"f3",X"22",X"f3",X"4e",X"8b",X"3c",X"0b",X"0b",X"3c",X"0b",X"0b",X"30",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"0d",X"f0",X"9e",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"b2",X"2e",X"54",X"62",X"51",X"62",X"cf",X"15",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"cf",X"62",X"15",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"51",X"62",X"51",X"61",X"2e",X"03",X"75",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"75",X"03",X"19",X"3c",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"12",X"aa",X"aa",X"98",X"83",X"0b",X"3c",X"2f",X"2e",X"1b",X"f0",X"6d",X"6d",X"aa",X"7c",X"aa",X"7c",X"9e",X"aa",X"a7",X"0c",X"a7",X"0b",X"d6",X"d6",X"32",X"e9",X"4d",X"e9",X"4d",X"bc",X"0b",X"0b",X"1b",X"0b",X"d1",X"4e",X"8b",X"d1",X"d1",X"57",X"82",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"54",X"ed",X"54",X"1b",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"3c",X"2f",X"54",X"3f",X"0b",X"1b",X"17",X"1b",X"00",X"0b",X"3c",X"0b",X"f3",X"ae",X"82",X"ae",X"ae",X"39",X"d1",X"d1",X"d1",X"d1",X"57",X"d1",X"d1",X"d1",X"0b",X"1b",X"0b",X"3c",X"0b",X"00",X"0b",X"eb",X"f3",X"f3",X"6f",X"af",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"2e",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"19",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"4f",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"3b",X"6d",X"f0",X"6d",X"6d",X"aa",X"aa",X"12",X"aa",X"98",X"0b",X"0b",X"0b",X"19",X"71",X"19",X"71",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"27",X"1a",X"03",X"03",X"1a",X"03",X"e5",X"2f",X"62",X"62",X"15",X"f5",X"51",X"62",X"51",X"cf",X"62",X"62",X"15",X"62",X"62",X"62",X"62",X"51",X"15",X"62",X"cf",X"62",X"15",X"cf",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"19",X"71",X"19",X"19",X"71",X"19",X"71",X"27",X"1a",X"03",X"19",X"03",X"19",X"b2",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"03",X"03",X"b2",X"ad",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",
    X"aa",X"2c",X"aa",X"60",X"61",X"0b",X"1b",X"83",X"69",X"ed",X"0b",X"6d",X"3f",X"f0",X"9e",X"aa",X"9e",X"aa",X"aa",X"7c",X"5f",X"36",X"0c",X"0b",X"2f",X"14",X"4d",X"e9",X"4d",X"bc",X"ea",X"0b",X"0b",X"e4",X"f3",X"d1",X"8b",X"39",X"1b",X"0b",X"65",X"6f",X"3c",X"54",X"2f",X"f0",X"0b",X"3c",X"2f",X"54",X"2f",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"0b",X"0b",X"00",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"54",X"2f",X"54",X"f0",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"00",X"0b",X"f3",X"ae",X"ae",X"39",X"ae",X"39",X"39",X"d1",X"d1",X"d1",X"57",X"39",X"d1",X"39",X"b8",X"0b",X"1b",X"0b",X"0b",X"0b",X"00",X"0b",X"3c",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"0b",X"3c",X"2e",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"f4",X"3c",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"92",X"aa",X"60",X"ba",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"75",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"2e",X"2f",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"51",X"f5",X"51",X"cf",X"15",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"f5",X"51",X"62",X"51",X"62",X"62",X"ed",X"2e",X"03",X"19",X"03",X"b2",X"03",X"19",X"71",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"75",X"03",X"1a",X"03",X"b2",X"19",X"3c",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"12",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"16",X"3c",X"98",X"f0",X"6d",X"6d",X"aa",X"7c",X"aa",X"1b",X"54",X"9e",X"a7",X"90",X"0c",X"3f",X"0b",X"ea",X"42",X"ea",X"fc",X"ea",X"54",X"1b",X"ae",X"82",X"82",X"57",X"d1",X"0b",X"d1",X"0b",X"1b",X"1b",X"54",X"2f",X"0b",X"54",X"2f",X"0b",X"54",X"f0",X"0b",X"00",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"00",X"1b",X"0b",X"0b",X"1b",X"3c",X"0b",X"3c",X"0b",X"3c",X"0b",X"3c",X"0b",X"3c",X"0b",X"2f",X"54",X"54",X"3f",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"3c",X"0b",X"f3",X"ae",X"82",X"39",X"39",X"fb",X"39",X"d1",X"57",X"d1",X"d1",X"39",X"d1",X"39",X"39",X"0b",X"0b",X"e4",X"1b",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"30",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"4a",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"3f",X"60",X"aa",X"aa",X"aa",X"98",X"1b",X"0b",X"0b",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"71",X"75",X"03",X"19",X"03",X"b2",X"d8",X"75",X"03",X"19",X"03",X"cc",X"54",X"62",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"f5",X"15",X"62",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"62",X"62",X"51",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"19",X"03",X"19",X"03",X"1a",X"03",X"b2",X"27",X"75",X"03",X"b2",X"d8",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"0b",X"0b",X"3c",X"33",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"7c",X"aa",X"ba",X"0b",X"1b",X"0b",X"69",X"0b",X"54",X"f0",X"6d",X"f0",X"aa",X"9e",X"0b",X"4d",X"1b",X"2f",X"a7",X"5f",X"68",X"36",X"0b",X"0b",X"1b",X"3c",X"0b",X"0b",X"3c",X"d6",X"0b",X"ae",X"ae",X"57",X"eb",X"39",X"d1",X"0b",X"d1",X"0b",X"f0",X"98",X"2f",X"0b",X"0b",X"54",X"2f",X"54",X"1b",X"0b",X"0b",X"00",X"0b",X"3c",X"0b",X"0b",X"0b",X"00",X"0b",X"1b",X"0b",X"54",X"98",X"54",X"2f",X"54",X"54",X"f0",X"0b",X"3c",X"0b",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"2f",X"2f",X"54",X"f0",X"0b",X"4e",X"af",X"6f",X"f3",X"f3",X"f3",X"ae",X"ae",X"39",X"ae",X"39",X"39",X"d1",X"d1",X"d1",X"d1",X"39",X"1f",X"39",X"4a",X"ae",X"39",X"ae",X"0b",X"0b",X"3c",X"0b",X"00",X"0b",X"3c",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"2e",X"03",X"1a",X"03",X"19",X"71",X"19",X"71",X"19",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"6d",X"aa",X"aa",X"7c",X"9e",X"98",X"0b",X"0b",X"0b",X"03",X"b2",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"75",X"03",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"2e",X"2f",X"62",X"51",X"62",X"cf",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"cf",X"62",X"62",X"15",X"cf",X"15",X"62",X"51",X"f0",X"2e",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"b2",X"27",X"19",X"71",X"19",X"03",X"19",X"03",X"03",X"b2",X"19",X"1b",X"0b",X"0b",X"53",X"6d",X"f0",X"3f",X"6d",
    X"aa",X"2c",X"aa",X"9e",X"54",X"0b",X"0b",X"0b",X"8c",X"0b",X"2f",X"6d",X"f0",X"6d",X"9e",X"aa",X"0b",X"fc",X"4d",X"0b",X"a7",X"36",X"0c",X"68",X"f0",X"a7",X"0c",X"2e",X"d6",X"f0",X"0b",X"d6",X"1b",X"0b",X"d1",X"0b",X"8b",X"ae",X"57",X"65",X"39",X"0b",X"54",X"2f",X"54",X"2f",X"0b",X"2f",X"98",X"2f",X"0b",X"0b",X"3c",X"0b",X"0b",X"0b",X"0b",X"3c",X"0b",X"1b",X"54",X"54",X"2f",X"f0",X"2f",X"f0",X"ed",X"54",X"2f",X"54",X"54",X"f0",X"0b",X"3c",X"0b",X"00",X"0b",X"0b",X"3c",X"0b",X"54",X"2f",X"6d",X"3c",X"0b",X"8b",X"f3",X"4e",X"f3",X"ae",X"f3",X"ae",X"ae",X"39",X"d1",X"4a",X"39",X"d1",X"ff",X"d1",X"57",X"39",X"d1",X"39",X"39",X"ae",X"82",X"ae",X"f3",X"0b",X"1b",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"0b",X"3c",X"2e",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"03",X"19",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"82",X"f4",X"91",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"3f",X"aa",X"60",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"71",X"19",X"03",X"19",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"cc",X"54",X"62",X"15",X"51",X"62",X"51",X"62",X"51",X"cf",X"62",X"62",X"62",X"15",X"f5",X"51",X"62",X"62",X"51",X"cf",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"0b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"12",X"aa",X"aa",X"84",X"0b",X"0b",X"1b",X"16",X"3c",X"98",X"f0",X"6d",X"f0",X"aa",X"7c",X"3c",X"0b",X"0b",X"1b",X"a7",X"5f",X"68",X"0c",X"d6",X"d6",X"2e",X"2e",X"2e",X"aa",X"0b",X"d6",X"d6",X"3c",X"0b",X"57",X"d1",X"0b",X"ae",X"39",X"6f",X"1b",X"2f",X"54",X"f0",X"0b",X"1b",X"54",X"f0",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"3c",X"0b",X"3c",X"54",X"ed",X"54",X"2f",X"f0",X"98",X"6d",X"6d",X"6d",X"f0",X"54",X"f0",X"ed",X"54",X"2f",X"54",X"1b",X"0b",X"0b",X"00",X"0b",X"0b",X"1b",X"54",X"2f",X"6d",X"1b",X"eb",X"8b",X"f3",X"f3",X"f3",X"ae",X"82",X"39",X"ae",X"39",X"39",X"d1",X"39",X"d1",X"d1",X"39",X"d1",X"39",X"fb",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"8b",X"1b",X"0b",X"3c",X"0b",X"00",X"0b",X"3c",X"2e",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"6d",X"aa",X"aa",X"60",X"aa",X"84",X"0b",X"1b",X"0b",X"75",X"71",X"19",X"71",X"19",X"19",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"19",X"2e",X"2f",X"62",X"62",X"62",X"15",X"62",X"62",X"62",X"62",X"15",X"cf",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"15",X"cf",X"15",X"f5",X"51",X"62",X"15",X"f5",X"62",X"15",X"cf",X"62",X"ed",X"2e",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"19",X"1b",X"0b",X"3c",X"17",X"f0",X"6d",X"3f",X"6d",
    X"aa",X"6d",X"aa",X"7c",X"61",X"0b",X"1b",X"83",X"69",X"0b",X"2f",X"6d",X"3f",X"6d",X"aa",X"9e",X"54",X"2f",X"aa",X"7c",X"9e",X"a7",X"36",X"0c",X"d6",X"d6",X"2e",X"2e",X"2e",X"0c",X"0b",X"d6",X"73",X"1b",X"0b",X"ae",X"82",X"d1",X"8b",X"1b",X"0b",X"00",X"d6",X"e9",X"2f",X"0b",X"2f",X"54",X"2f",X"0b",X"00",X"0b",X"3c",X"0b",X"3c",X"0b",X"1b",X"54",X"f0",X"54",X"f0",X"6d",X"6d",X"6d",X"aa",X"aa",X"9e",X"1a",X"6d",X"f0",X"54",X"f0",X"54",X"2f",X"54",X"3c",X"0b",X"3c",X"0b",X"3c",X"0b",X"ed",X"54",X"f0",X"0b",X"0b",X"8b",X"4e",X"f3",X"ae",X"f3",X"ae",X"ae",X"39",X"fb",X"39",X"d1",X"d1",X"57",X"d1",X"57",X"4a",X"57",X"39",X"39",X"ae",X"82",X"ae",X"f3",X"f3",X"22",X"f3",X"4e",X"0b",X"1b",X"0b",X"0b",X"00",X"0b",X"2e",X"19",X"03",X"b2",X"03",X"75",X"03",X"03",X"1a",X"03",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"9e",X"7c",X"aa",X"aa",X"98",X"0b",X"0b",X"0b",X"03",X"03",X"19",X"03",X"b2",X"27",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"75",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"2e",X"ed",X"51",X"62",X"51",X"62",X"cf",X"15",X"51",X"f5",X"51",X"62",X"15",X"f5",X"51",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"77",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"b2",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"0b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"36",X"9e",X"aa",X"98",X"0b",X"0b",X"1b",X"16",X"1b",X"98",X"f0",X"6d",X"f0",X"6d",X"aa",X"92",X"aa",X"6d",X"aa",X"aa",X"a7",X"a7",X"89",X"d6",X"d6",X"2e",X"2e",X"ec",X"d6",X"0b",X"ea",X"0b",X"0b",X"ae",X"70",X"ff",X"f3",X"0b",X"d1",X"ff",X"0b",X"2e",X"2e",X"4d",X"1b",X"54",X"2f",X"54",X"1b",X"0b",X"0b",X"0b",X"0b",X"3c",X"0b",X"ed",X"54",X"2f",X"6d",X"1a",X"6d",X"9e",X"aa",X"aa",X"60",X"aa",X"92",X"aa",X"6d",X"6d",X"f0",X"98",X"f0",X"54",X"f0",X"0b",X"0b",X"0b",X"3c",X"0b",X"3c",X"54",X"54",X"f0",X"0b",X"af",X"f3",X"4e",X"f3",X"ae",X"ae",X"39",X"ae",X"39",X"39",X"d1",X"d1",X"d1",X"d1",X"d1",X"ff",X"39",X"4a",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"f3",X"f3",X"6f",X"af",X"8b",X"0b",X"3c",X"0b",X"0b",X"3c",X"2e",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"9e",X"aa",X"9e",X"98",X"0b",X"0b",X"3c",X"03",X"19",X"b2",X"27",X"19",X"b2",X"03",X"1a",X"03",X"03",X"19",X"b2",X"03",X"03",X"1a",X"71",X"19",X"71",X"27",X"1a",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"ec",X"f0",X"62",X"62",X"62",X"62",X"51",X"62",X"15",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"cf",X"62",X"15",X"51",X"62",X"62",X"15",X"61",X"2e",X"1a",X"03",X"19",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"1b",X"0b",X"1b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"60",X"aa",X"60",X"98",X"1b",X"1b",X"0b",X"69",X"00",X"54",X"f0",X"6d",X"3f",X"54",X"aa",X"aa",X"9e",X"36",X"9e",X"6d",X"a7",X"5f",X"68",X"0c",X"d6",X"d6",X"2e",X"2e",X"2e",X"3c",X"0b",X"ae",X"82",X"ae",X"82",X"ae",X"57",X"57",X"39",X"d1",X"0b",X"2f",X"42",X"d6",X"0b",X"f0",X"98",X"0b",X"00",X"0b",X"3c",X"0b",X"00",X"0b",X"54",X"f0",X"2f",X"6d",X"3f",X"6d",X"aa",X"aa",X"a7",X"6d",X"a7",X"aa",X"36",X"9e",X"aa",X"aa",X"6d",X"f0",X"6d",X"2f",X"54",X"2f",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"2f",X"54",X"3f",X"0b",X"8b",X"f3",X"f3",X"f3",X"ae",X"70",X"39",X"39",X"fb",X"39",X"d1",X"d1",X"57",X"d1",X"39",X"d1",X"d1",X"39",X"ae",X"82",X"b7",X"f3",X"f3",X"46",X"8b",X"f3",X"4e",X"8b",X"3c",X"0b",X"0b",X"3c",X"0b",X"3c",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"7c",X"aa",X"7c",X"61",X"0b",X"1b",X"0b",X"75",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"2e",X"54",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"cf",X"62",X"62",X"62",X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"cf",X"62",X"62",X"51",X"62",X"77",X"2e",X"03",X"03",X"b2",X"03",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"03",X"1a",X"03",X"19",X"03",X"06",X"03",X"1a",X"03",X"1a",X"03",X"0b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"aa",X"aa",X"aa",X"98",X"0b",X"0b",X"0b",X"79",X"2e",X"0b",X"f0",X"6d",X"f0",X"6d",X"9e",X"7c",X"aa",X"6d",X"aa",X"aa",X"a7",X"5f",X"68",X"0c",X"f8",X"d6",X"2e",X"2e",X"2e",X"1b",X"0b",X"3c",X"0b",X"ae",X"82",X"ae",X"82",X"ae",X"39",X"d1",X"8b",X"3c",X"98",X"ea",X"0b",X"2f",X"54",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"2f",X"54",X"6d",X"f0",X"6d",X"aa",X"9e",X"a7",X"6d",X"a7",X"3f",X"36",X"12",X"a7",X"aa",X"60",X"aa",X"6d",X"f0",X"98",X"f0",X"54",X"3c",X"0b",X"0b",X"3c",X"0b",X"3c",X"54",X"2f",X"6d",X"3c",X"f3",X"6f",X"f3",X"ae",X"f3",X"ae",X"ae",X"39",X"39",X"39",X"4a",X"57",X"d1",X"57",X"d1",X"39",X"4a",X"39",X"4a",X"ae",X"82",X"ae",X"f3",X"f3",X"f3",X"4e",X"8b",X"4e",X"0b",X"00",X"3c",X"0b",X"0b",X"3c",X"2e",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"91",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"cd",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"9e",X"aa",X"84",X"0b",X"0b",X"0b",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"03",X"2e",X"2f",X"62",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"41",X"8e",X"8e",X"b1",X"8e",X"8e",X"2d",X"41",X"51",X"62",X"62",X"15",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"ed",X"2e",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"03",X"1a",X"03",X"b2",X"27",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"03",X"1a",X"e4",X"0b",X"0b",X"3b",X"f0",X"6d",X"3f",X"6d",
    X"9e",X"7c",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"79",X"2e",X"1b",X"54",X"f0",X"6d",X"3f",X"aa",X"aa",X"aa",X"12",X"aa",X"7c",X"5f",X"a7",X"36",X"a7",X"aa",X"54",X"3c",X"1b",X"3c",X"0b",X"1b",X"d6",X"0b",X"3c",X"0b",X"8b",X"ae",X"82",X"39",X"fb",X"57",X"0b",X"3c",X"54",X"1b",X"54",X"2f",X"0b",X"0b",X"3c",X"0b",X"00",X"0b",X"2f",X"54",X"ed",X"f0",X"6d",X"aa",X"aa",X"90",X"aa",X"a7",X"5f",X"a7",X"90",X"5f",X"6d",X"a7",X"aa",X"9e",X"6d",X"f0",X"6d",X"2f",X"98",X"f0",X"0b",X"3c",X"0b",X"0b",X"0b",X"1b",X"54",X"f0",X"0b",X"4e",X"f3",X"f3",X"22",X"ae",X"ae",X"39",X"ae",X"d1",X"4a",X"57",X"39",X"d1",X"d1",X"39",X"d1",X"d1",X"39",X"ae",X"39",X"ae",X"f3",X"ae",X"f3",X"f3",X"22",X"8b",X"af",X"0b",X"0b",X"0b",X"0b",X"3c",X"0b",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"75",X"03",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"33",X"6d",X"3f",X"6d",X"f0",X"60",X"aa",X"7c",X"aa",X"98",X"0b",X"0b",X"1b",X"03",X"1a",X"b2",X"19",X"03",X"1a",X"03",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"03",X"75",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"2e",X"ed",X"62",X"51",X"62",X"cf",X"15",X"f5",X"15",X"62",X"62",X"15",X"62",X"41",X"8e",X"c7",X"8f",X"30",X"5b",X"18",X"41",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"79",X"2e",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"75",X"03",X"b2",X"03",X"1a",X"03",X"71",X"19",X"b2",X"03",X"19",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"06",X"19",X"b2",X"03",X"b2",X"19",X"1b",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"1b",X"83",X"2f",X"2e",X"0b",X"3c",X"6d",X"f0",X"6d",X"aa",X"9e",X"2c",X"f0",X"54",X"2f",X"0b",X"0b",X"3c",X"1b",X"0b",X"0b",X"0b",X"4d",X"e9",X"d6",X"d6",X"2e",X"d6",X"1b",X"3c",X"ae",X"82",X"ae",X"39",X"39",X"d1",X"ae",X"0b",X"1b",X"0b",X"2f",X"54",X"00",X"0b",X"0b",X"3c",X"0b",X"0b",X"2f",X"54",X"f0",X"6d",X"3f",X"6d",X"12",X"aa",X"a7",X"5f",X"90",X"a7",X"5f",X"5f",X"a7",X"6d",X"aa",X"7c",X"9e",X"1a",X"6d",X"54",X"2f",X"54",X"1b",X"0b",X"3c",X"0b",X"00",X"0b",X"2f",X"54",X"0b",X"f3",X"8b",X"f3",X"ae",X"f3",X"ae",X"82",X"39",X"39",X"39",X"fb",X"d1",X"ff",X"d1",X"57",X"39",X"4a",X"39",X"39",X"ae",X"ae",X"82",X"f3",X"f3",X"22",X"48",X"f3",X"4e",X"8b",X"1b",X"0b",X"00",X"0b",X"0b",X"2e",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"9e",X"aa",X"84",X"0b",X"0b",X"1b",X"19",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"19",X"b2",X"27",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"2e",X"2f",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"cf",X"62",X"41",X"8e",X"a4",X"30",X"18",X"30",X"8e",X"41",X"51",X"62",X"15",X"cf",X"62",X"15",X"51",X"62",X"62",X"51",X"62",X"62",X"ed",X"2e",X"03",X"03",X"19",X"03",X"03",X"b2",X"27",X"19",X"71",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"03",X"03",X"b2",X"27",X"75",X"03",X"03",X"03",X"03",X"03",X"19",X"03",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"12",X"98",X"0b",X"0b",X"1b",X"ed",X"03",X"2e",X"3c",X"6d",X"f0",X"6d",X"3c",X"0b",X"3c",X"1b",X"0b",X"00",X"1b",X"0b",X"0b",X"0b",X"0b",X"1b",X"3c",X"0b",X"aa",X"d6",X"d6",X"d6",X"d6",X"ad",X"8b",X"ae",X"70",X"ae",X"82",X"d1",X"39",X"d1",X"d1",X"8b",X"3c",X"54",X"2f",X"0b",X"0b",X"3c",X"0b",X"0b",X"1b",X"54",X"2f",X"54",X"f0",X"6d",X"aa",X"aa",X"a7",X"3f",X"a7",X"36",X"5f",X"a7",X"90",X"aa",X"a7",X"9e",X"aa",X"aa",X"6d",X"3f",X"2f",X"54",X"54",X"1b",X"0b",X"0b",X"3c",X"0b",X"0b",X"ed",X"54",X"1b",X"4e",X"f3",X"f3",X"f3",X"ae",X"70",X"d1",X"ae",X"39",X"4a",X"57",X"39",X"d1",X"d1",X"d1",X"d1",X"39",X"d1",X"82",X"39",X"ae",X"f3",X"ae",X"f3",X"f3",X"f3",X"6f",X"8b",X"af",X"0b",X"1b",X"0b",X"0b",X"3c",X"0b",X"ec",X"03",X"b2",X"03",X"03",X"03",X"19",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"70",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",X"12",X"aa",X"7c",X"aa",X"98",X"1b",X"0b",X"0b",X"d8",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"2e",X"54",X"62",X"51",X"15",X"62",X"15",X"51",X"62",X"62",X"62",X"15",X"f5",X"f5",X"8e",X"30",X"5b",X"c7",X"8f",X"18",X"41",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"f5",X"51",X"f0",X"2e",X"03",X"19",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"75",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"19",X"b2",X"19",X"b2",X"d8",X"0b",X"1b",X"0b",X"33",X"6d",X"f0",X"3f",X"6d",
    X"9e",X"aa",X"9e",X"aa",X"98",X"0b",X"1b",X"0b",X"2f",X"03",X"cc",X"0b",X"1b",X"0b",X"3c",X"0b",X"1b",X"0b",X"0b",X"0b",X"54",X"6d",X"aa",X"0c",X"0c",X"f8",X"d6",X"68",X"aa",X"0b",X"0b",X"d6",X"4d",X"1b",X"82",X"ae",X"82",X"ae",X"b7",X"ae",X"82",X"39",X"39",X"d1",X"d1",X"0b",X"1b",X"54",X"f0",X"0b",X"3c",X"0b",X"2f",X"54",X"f0",X"54",X"54",X"f0",X"6d",X"aa",X"7c",X"6d",X"a7",X"90",X"5f",X"a7",X"36",X"a7",X"5f",X"aa",X"2c",X"aa",X"9e",X"6d",X"f0",X"54",X"f0",X"58",X"3c",X"0b",X"0b",X"3c",X"0b",X"1b",X"54",X"2f",X"0b",X"f3",X"6f",X"22",X"ae",X"f3",X"ae",X"82",X"39",X"39",X"d1",X"39",X"d1",X"ff",X"d1",X"d1",X"39",X"39",X"4a",X"39",X"ae",X"82",X"ae",X"f3",X"f3",X"22",X"8b",X"e0",X"4e",X"8b",X"3c",X"0b",X"00",X"0b",X"00",X"0b",X"2e",X"1a",X"03",X"03",X"b2",X"19",X"b2",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"60",X"aa",X"92",X"61",X"0b",X"0b",X"1b",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"ec",X"2f",X"62",X"62",X"62",X"62",X"cf",X"62",X"62",X"51",X"62",X"51",X"62",X"f5",X"18",X"5b",X"18",X"30",X"c7",X"18",X"34",X"15",X"f5",X"62",X"51",X"62",X"cf",X"62",X"15",X"51",X"62",X"62",X"15",X"61",X"2e",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"03",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"f0",X"6d",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"79",X"03",X"19",X"ec",X"0b",X"3c",X"2e",X"2e",X"3c",X"54",X"f0",X"aa",X"9e",X"aa",X"5f",X"a7",X"89",X"0c",X"d6",X"d6",X"2e",X"0c",X"aa",X"0b",X"e9",X"3c",X"3c",X"0b",X"82",X"ae",X"82",X"70",X"ae",X"d1",X"4a",X"39",X"d1",X"ae",X"0b",X"54",X"2f",X"0b",X"0b",X"fc",X"d6",X"2e",X"d6",X"fc",X"2f",X"98",X"2f",X"9e",X"aa",X"5f",X"aa",X"a7",X"5f",X"90",X"5f",X"a7",X"6d",X"a7",X"9e",X"aa",X"6d",X"f0",X"6d",X"ed",X"54",X"f0",X"0b",X"00",X"3c",X"0b",X"0b",X"3c",X"54",X"f0",X"0b",X"af",X"f3",X"f3",X"f3",X"ae",X"ae",X"39",X"ae",X"39",X"4a",X"d1",X"39",X"57",X"d1",X"39",X"d1",X"d1",X"0b",X"3c",X"0b",X"0b",X"0b",X"eb",X"8b",X"f3",X"f3",X"8b",X"8b",X"8b",X"3c",X"1b",X"0b",X"0b",X"0b",X"1b",X"2e",X"03",X"03",X"1a",X"03",X"03",X"03",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"91",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"2e",X"54",X"62",X"51",X"62",X"51",X"62",X"15",X"cf",X"62",X"15",X"62",X"62",X"f5",X"24",X"18",X"30",X"24",X"18",X"18",X"41",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"ed",X"2e",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"71",X"19",X"b2",X"27",X"19",X"03",X"19",X"03",X"b2",X"d8",X"19",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"19",X"b2",X"19",X"0b",X"1b",X"0b",X"53",X"6d",X"f0",X"3f",X"6d",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"77",X"03",X"b2",X"2e",X"2e",X"2e",X"1b",X"0b",X"2f",X"60",X"aa",X"7c",X"aa",X"7c",X"aa",X"a7",X"0c",X"0c",X"f8",X"d6",X"2e",X"2e",X"d6",X"aa",X"14",X"4d",X"bc",X"0b",X"3c",X"1b",X"82",X"ae",X"82",X"39",X"39",X"39",X"fb",X"57",X"0b",X"2f",X"54",X"3c",X"0b",X"d6",X"2e",X"ec",X"2e",X"2e",X"d6",X"fc",X"54",X"f0",X"9e",X"36",X"90",X"aa",X"a7",X"aa",X"a7",X"9e",X"a7",X"aa",X"aa",X"7c",X"f0",X"6d",X"f0",X"54",X"2f",X"54",X"1b",X"0b",X"0b",X"0b",X"3c",X"0b",X"54",X"2f",X"0b",X"0b",X"eb",X"f3",X"ae",X"f3",X"ae",X"ae",X"39",X"d1",X"39",X"39",X"d1",X"d1",X"d1",X"57",X"4a",X"39",X"f3",X"0b",X"1b",X"3c",X"0b",X"3c",X"0b",X"0b",X"3c",X"eb",X"4e",X"eb",X"0b",X"0b",X"3c",X"0b",X"3c",X"2e",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"cd",X"6d",X"3f",X"98",X"6d",X"aa",X"12",X"6d",X"12",X"98",X"0b",X"0b",X"0b",X"19",X"71",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"03",X"19",X"b2",X"27",X"19",X"03",X"b2",X"03",X"e5",X"2f",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"0f",X"18",X"5b",X"5b",X"18",X"5b",X"8e",X"f5",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"15",X"cf",X"62",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"03",X"75",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"71",X"03",X"19",X"b2",X"27",X"19",X"b2",X"27",X"19",X"03",X"03",X"b2",X"19",X"03",X"03",X"03",X"0b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"0d",X"60",X"61",X"0b",X"0b",X"0b",X"2f",X"03",X"1a",X"2e",X"1b",X"0b",X"54",X"3f",X"6d",X"aa",X"aa",X"9e",X"aa",X"9e",X"aa",X"90",X"5f",X"89",X"0c",X"f8",X"d6",X"2e",X"2e",X"0c",X"1b",X"42",X"ea",X"fc",X"0b",X"8b",X"ae",X"82",X"b7",X"82",X"39",X"d1",X"39",X"d1",X"ae",X"0b",X"f0",X"54",X"1b",X"f8",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"f0",X"6d",X"aa",X"9e",X"aa",X"a7",X"6d",X"a7",X"aa",X"a7",X"6d",X"aa",X"12",X"f0",X"6d",X"3f",X"54",X"f0",X"54",X"2f",X"0b",X"0b",X"3c",X"00",X"0b",X"3c",X"ed",X"54",X"1b",X"0b",X"0b",X"af",X"f3",X"ae",X"82",X"39",X"ae",X"39",X"4a",X"d1",X"d1",X"d1",X"57",X"d1",X"57",X"39",X"4a",X"39",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"00",X"0b",X"0b",X"0b",X"00",X"0b",X"3c",X"0b",X"30",X"03",X"03",X"19",X"03",X"71",X"19",X"03",X"19",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"60",X"aa",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"1a",X"03",X"03",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"75",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"2e",X"ed",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"51",X"62",X"cf",X"62",X"a1",X"18",X"5b",X"18",X"18",X"5b",X"18",X"0f",X"62",X"51",X"cf",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"79",X"2e",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"71",X"19",X"b2",X"1b",X"0b",X"0b",X"17",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"7c",X"aa",X"84",X"0b",X"0b",X"1b",X"61",X"03",X"03",X"2e",X"3c",X"f0",X"3f",X"6d",X"f0",X"9e",X"7c",X"aa",X"7c",X"aa",X"9e",X"a7",X"5f",X"a7",X"0c",X"0c",X"d6",X"d6",X"2e",X"2e",X"aa",X"6d",X"fc",X"ea",X"0b",X"ae",X"82",X"ae",X"82",X"ae",X"82",X"ae",X"39",X"39",X"d1",X"82",X"0b",X"2f",X"0b",X"3c",X"2e",X"2e",X"2e",X"ec",X"2e",X"2e",X"d6",X"6d",X"f0",X"6d",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"9e",X"f0",X"6d",X"6d",X"f0",X"6d",X"2f",X"54",X"2f",X"0b",X"0b",X"3c",X"0b",X"0b",X"0b",X"54",X"f0",X"6d",X"00",X"2e",X"00",X"0b",X"eb",X"f3",X"ae",X"ae",X"39",X"39",X"d1",X"39",X"d1",X"ff",X"d1",X"57",X"4a",X"d1",X"39",X"d1",X"4a",X"ae",X"0b",X"e4",X"0b",X"1b",X"0b",X"0b",X"3c",X"1b",X"0b",X"0b",X"2e",X"2e",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"7c",X"9e",X"98",X"0b",X"0b",X"3c",X"d8",X"75",X"03",X"03",X"71",X"19",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"75",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"27",X"2e",X"2f",X"62",X"15",X"62",X"cf",X"62",X"62",X"62",X"62",X"15",X"62",X"62",X"f5",X"8e",X"24",X"18",X"24",X"18",X"8e",X"0f",X"62",X"62",X"62",X"15",X"62",X"62",X"51",X"15",X"62",X"62",X"15",X"62",X"ed",X"2e",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"71",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"0b",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"2f",X"03",X"1a",X"ec",X"0b",X"54",X"6d",X"f0",X"6d",X"f0",X"aa",X"60",X"aa",X"aa",X"7c",X"aa",X"a7",X"5f",X"68",X"0c",X"d6",X"d6",X"2e",X"2e",X"0c",X"0b",X"ea",X"fc",X"0b",X"82",X"6f",X"3c",X"0b",X"8b",X"ae",X"70",X"ae",X"d1",X"d1",X"57",X"0b",X"54",X"0b",X"1b",X"42",X"d6",X"2e",X"2e",X"2e",X"2e",X"d6",X"2f",X"6d",X"f0",X"6d",X"3f",X"aa",X"9e",X"aa",X"6d",X"f0",X"6d",X"f0",X"f0",X"98",X"2f",X"54",X"2f",X"54",X"0b",X"00",X"0b",X"0b",X"1b",X"0b",X"2f",X"54",X"f0",X"0b",X"2e",X"2e",X"0b",X"3c",X"0b",X"82",X"39",X"ae",X"39",X"4a",X"39",X"39",X"d1",X"d1",X"d1",X"ff",X"39",X"fb",X"39",X"ae",X"39",X"ae",X"82",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"2e",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"70",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"c6",X"6d",X"f0",X"3f",X"6d",X"aa",X"9e",X"aa",X"aa",X"74",X"0b",X"0b",X"1b",X"19",X"71",X"27",X"19",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"b2",X"27",X"19",X"03",X"b2",X"2e",X"98",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"51",X"62",X"51",X"62",X"a1",X"18",X"18",X"24",X"18",X"18",X"8e",X"f5",X"51",X"62",X"51",X"62",X"cf",X"15",X"62",X"62",X"62",X"51",X"62",X"51",X"f0",X"2e",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"19",X"03",X"03",X"b2",X"03",X"19",X"71",X"03",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"19",X"b2",X"27",X"19",X"03",X"b2",X"19",X"1b",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",
    X"aa",X"7c",X"aa",X"9e",X"98",X"0b",X"0b",X"0b",X"77",X"03",X"19",X"71",X"2e",X"1b",X"f0",X"6d",X"6d",X"f0",X"12",X"aa",X"aa",X"9e",X"54",X"2f",X"0b",X"54",X"5f",X"0c",X"68",X"d6",X"d6",X"2e",X"2e",X"1b",X"9e",X"36",X"1b",X"3c",X"1b",X"0b",X"3c",X"ae",X"82",X"ae",X"82",X"70",X"d1",X"d1",X"ae",X"0b",X"2f",X"0b",X"0b",X"3c",X"42",X"d6",X"2e",X"d6",X"42",X"f0",X"54",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"3f",X"54",X"54",X"f0",X"54",X"f0",X"54",X"3c",X"1b",X"0b",X"0b",X"00",X"0b",X"2f",X"54",X"ed",X"6d",X"1b",X"2e",X"03",X"21",X"1b",X"0b",X"3c",X"82",X"39",X"d1",X"39",X"4a",X"d1",X"39",X"ff",X"d1",X"39",X"d1",X"39",X"39",X"39",X"ae",X"ae",X"ae",X"f3",X"0b",X"1b",X"0b",X"3c",X"0b",X"0b",X"00",X"0b",X"0b",X"3c",X"2e",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"91",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"7c",X"9e",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"19",X"71",X"19",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"03",X"19",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"ec",X"2f",X"51",X"62",X"62",X"15",X"f5",X"51",X"62",X"62",X"62",X"62",X"62",X"51",X"18",X"ff",X"18",X"f9",X"8e",X"8e",X"a1",X"62",X"62",X"62",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"62",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"1a",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"0b",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"9e",X"2c",X"ba",X"0b",X"1b",X"83",X"2f",X"03",X"b2",X"19",X"2e",X"00",X"6d",X"3f",X"f0",X"6d",X"f0",X"2f",X"0b",X"0b",X"21",X"2e",X"2e",X"1b",X"aa",X"68",X"0c",X"f8",X"d6",X"2e",X"2e",X"0b",X"aa",X"fc",X"d6",X"2e",X"2e",X"2e",X"1b",X"82",X"ae",X"ae",X"82",X"ae",X"ae",X"39",X"d1",X"ae",X"54",X"2f",X"0b",X"0b",X"3c",X"2f",X"54",X"2f",X"0b",X"ed",X"54",X"2f",X"54",X"6d",X"f0",X"6d",X"f0",X"6d",X"f0",X"54",X"2f",X"54",X"2f",X"54",X"ed",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"54",X"f0",X"6d",X"3c",X"2e",X"03",X"19",X"03",X"2e",X"3c",X"0b",X"3c",X"82",X"39",X"4f",X"39",X"d1",X"d1",X"d1",X"d1",X"ff",X"39",X"fb",X"39",X"ae",X"39",X"ae",X"70",X"ae",X"f3",X"f3",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"2e",X"03",X"19",X"03",X"1a",X"03",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"9e",X"aa",X"7c",X"53",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"03",X"2e",X"98",X"62",X"62",X"51",X"62",X"15",X"62",X"cf",X"0f",X"a1",X"a1",X"0f",X"34",X"18",X"8e",X"18",X"8e",X"18",X"8e",X"51",X"a1",X"f5",X"a1",X"51",X"62",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"ed",X"2e",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"d8",X"0b",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"ed",X"03",X"19",X"03",X"2e",X"1b",X"54",X"f0",X"6d",X"ed",X"0b",X"6d",X"30",X"2e",X"03",X"03",X"cc",X"0b",X"a7",X"36",X"0c",X"0c",X"f8",X"d6",X"2e",X"3c",X"aa",X"2e",X"2e",X"2e",X"ec",X"e9",X"3c",X"ae",X"8b",X"3c",X"0b",X"ae",X"82",X"8b",X"1b",X"0b",X"3c",X"98",X"2f",X"0b",X"0b",X"0b",X"0b",X"00",X"0b",X"3c",X"0b",X"ed",X"54",X"2f",X"54",X"f0",X"54",X"2f",X"54",X"2f",X"54",X"2f",X"54",X"1b",X"0b",X"3c",X"0b",X"3c",X"0b",X"3c",X"0b",X"54",X"2f",X"54",X"f0",X"0b",X"21",X"03",X"b2",X"03",X"1a",X"2e",X"3c",X"0b",X"0b",X"af",X"39",X"39",X"d1",X"39",X"d1",X"57",X"39",X"d1",X"39",X"39",X"d1",X"82",X"ae",X"ae",X"f3",X"ae",X"f3",X"f3",X"1b",X"0b",X"3c",X"0b",X"00",X"0b",X"0b",X"3c",X"0b",X"0b",X"30",X"03",X"b2",X"03",X"03",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"70",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",X"7c",X"aa",X"aa",X"12",X"98",X"0b",X"1b",X"0b",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"75",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"d8",X"19",X"71",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"03",X"b2",X"2e",X"2f",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"51",X"18",X"8e",X"8e",X"8e",X"18",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"41",X"a1",X"51",X"62",X"51",X"62",X"cf",X"15",X"62",X"15",X"54",X"2e",X"19",X"71",X"27",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"71",X"19",X"b2",X"27",X"19",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"b2",X"cd",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",
    X"aa",X"9e",X"aa",X"9e",X"98",X"1b",X"0b",X"0b",X"2f",X"03",X"b2",X"03",X"b2",X"2e",X"1b",X"0b",X"1b",X"6d",X"2e",X"ec",X"03",X"03",X"cc",X"2e",X"0b",X"aa",X"90",X"5f",X"68",X"0c",X"d6",X"d6",X"f8",X"0b",X"2e",X"2e",X"2e",X"ec",X"73",X"2f",X"0b",X"1b",X"1b",X"d6",X"3c",X"f3",X"0b",X"0b",X"1b",X"b8",X"f3",X"0b",X"f0",X"54",X"3c",X"0b",X"3c",X"0b",X"0b",X"0b",X"3c",X"0b",X"3c",X"54",X"2f",X"54",X"2f",X"54",X"2f",X"54",X"1b",X"0b",X"3c",X"0b",X"0b",X"0b",X"3c",X"0b",X"0b",X"0b",X"f0",X"2f",X"54",X"f0",X"0b",X"2e",X"03",X"19",X"03",X"1a",X"03",X"03",X"cc",X"fc",X"1b",X"0b",X"65",X"39",X"d1",X"d1",X"d1",X"d1",X"d1",X"d1",X"39",X"fb",X"82",X"39",X"ae",X"82",X"ae",X"f3",X"f3",X"f3",X"6f",X"f3",X"0b",X"1b",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"2e",X"03",X"1a",X"03",X"1a",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"9e",X"aa",X"2c",X"aa",X"61",X"0b",X"0b",X"0b",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"71",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"2e",X"ed",X"62",X"62",X"15",X"62",X"62",X"15",X"51",X"62",X"51",X"18",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"41",X"a1",X"62",X"62",X"15",X"f5",X"62",X"51",X"62",X"cf",X"62",X"f0",X"2e",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"71",X"19",X"03",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"27",X"27",X"0b",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"7c",X"61",X"0b",X"0b",X"1b",X"61",X"03",X"75",X"03",X"19",X"2e",X"3c",X"54",X"2e",X"ec",X"03",X"19",X"2e",X"2e",X"3c",X"0b",X"aa",X"9e",X"aa",X"a7",X"5f",X"68",X"0c",X"d6",X"0c",X"e4",X"2e",X"2e",X"4d",X"f0",X"54",X"fc",X"d6",X"32",X"e9",X"4d",X"1b",X"0b",X"3c",X"eb",X"f3",X"8b",X"46",X"f3",X"0b",X"ed",X"54",X"2f",X"0b",X"1b",X"0b",X"00",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"0b",X"0b",X"00",X"0b",X"3c",X"0b",X"0b",X"00",X"0b",X"00",X"0b",X"0b",X"3c",X"2f",X"54",X"98",X"f0",X"6d",X"0b",X"30",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"b2",X"2e",X"3c",X"0b",X"3c",X"d1",X"39",X"ff",X"d1",X"39",X"d1",X"39",X"39",X"4a",X"ae",X"82",X"b7",X"f3",X"ae",X"f3",X"22",X"f3",X"af",X"8b",X"4e",X"0b",X"0b",X"00",X"0b",X"0b",X"3c",X"0b",X"ec",X"03",X"03",X"03",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"84",X"f0",X"6d",X"3f",X"6d",X"aa",X"9e",X"aa",X"7c",X"33",X"0b",X"1b",X"0b",X"d8",X"1a",X"03",X"03",X"b2",X"27",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"71",X"19",X"b2",X"03",X"27",X"19",X"71",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"75",X"03",X"03",X"b2",X"03",X"19",X"2e",X"2f",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"51",X"18",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"51",X"15",X"62",X"cf",X"62",X"51",X"15",X"62",X"62",X"62",X"51",X"2f",X"2e",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"19",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"1b",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"9e",X"aa",X"98",X"0b",X"1b",X"0b",X"2f",X"03",X"b2",X"03",X"b2",X"03",X"e5",X"2e",X"03",X"1a",X"2e",X"ec",X"0b",X"1b",X"9e",X"aa",X"7c",X"aa",X"9e",X"a7",X"36",X"68",X"0c",X"68",X"1b",X"0b",X"4d",X"f0",X"54",X"fc",X"d6",X"d6",X"d6",X"73",X"4d",X"fc",X"1b",X"0b",X"4e",X"8b",X"4e",X"f3",X"f3",X"f3",X"f3",X"ad",X"1b",X"54",X"54",X"3c",X"1b",X"0b",X"0b",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"1b",X"0b",X"00",X"0b",X"0b",X"00",X"0b",X"1b",X"0b",X"0b",X"3c",X"54",X"54",X"2f",X"2f",X"6d",X"3c",X"cc",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"19",X"2e",X"3c",X"0b",X"0b",X"d1",X"d1",X"d1",X"ff",X"39",X"fb",X"39",X"d1",X"39",X"ae",X"82",X"ae",X"f3",X"82",X"f3",X"8b",X"22",X"8b",X"af",X"0b",X"1b",X"0b",X"0b",X"00",X"0b",X"0b",X"2e",X"19",X"b2",X"19",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"91",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"3b",X"6d",X"f0",X"6d",X"f0",X"7c",X"aa",X"9e",X"aa",X"98",X"0b",X"0b",X"0b",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"03",X"1a",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"30",X"f0",X"62",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"15",X"62",X"51",X"18",X"8e",X"8e",X"8e",X"8e",X"8e",X"8e",X"41",X"51",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"61",X"2e",X"03",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"19",X"0b",X"0b",X"0b",X"33",X"6d",X"3f",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"79",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"2e",X"2e",X"3c",X"0b",X"6d",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"aa",X"a7",X"5f",X"0c",X"0c",X"1b",X"42",X"f0",X"42",X"0b",X"d6",X"d6",X"14",X"4d",X"fc",X"42",X"3c",X"0b",X"0b",X"af",X"8b",X"f3",X"4e",X"f3",X"f3",X"ae",X"f3",X"ae",X"0b",X"2f",X"54",X"54",X"1b",X"0b",X"3c",X"3c",X"0b",X"00",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"1b",X"0b",X"0b",X"3c",X"0b",X"54",X"f0",X"ed",X"54",X"6d",X"00",X"2e",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"d8",X"30",X"1b",X"0b",X"1b",X"0b",X"d1",X"39",X"d1",X"39",X"4a",X"39",X"ae",X"39",X"ae",X"82",X"82",X"f3",X"f3",X"22",X"af",X"8b",X"4e",X"8b",X"00",X"0b",X"1b",X"0b",X"0b",X"3c",X"0b",X"2e",X"03",X"03",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",X"12",X"aa",X"7c",X"aa",X"84",X"0b",X"0b",X"3c",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"2e",X"54",X"51",X"62",X"15",X"62",X"15",X"f5",X"15",X"62",X"cf",X"62",X"51",X"51",X"18",X"8e",X"8e",X"8e",X"8e",X"5c",X"51",X"62",X"62",X"51",X"62",X"15",X"f5",X"15",X"cf",X"62",X"62",X"15",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"19",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"75",X"03",X"75",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"ed",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"2e",X"3c",X"0b",X"3f",X"6d",X"f0",X"9e",X"aa",X"aa",X"7c",X"aa",X"60",X"aa",X"12",X"36",X"0b",X"0b",X"4d",X"d6",X"2e",X"0c",X"aa",X"0b",X"0b",X"fc",X"42",X"bc",X"ea",X"0b",X"1b",X"65",X"8b",X"6f",X"af",X"f3",X"f3",X"22",X"f3",X"ae",X"82",X"b7",X"0b",X"0b",X"ed",X"54",X"2f",X"54",X"54",X"1b",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"0b",X"3c",X"54",X"2f",X"98",X"2f",X"54",X"2f",X"6d",X"3c",X"1b",X"cc",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"19",X"b2",X"27",X"2e",X"2e",X"00",X"0b",X"0b",X"3c",X"39",X"d1",X"39",X"4a",X"39",X"ae",X"82",X"b7",X"f3",X"ae",X"f3",X"f3",X"f3",X"6f",X"af",X"8b",X"1b",X"0b",X"00",X"0b",X"3c",X"0b",X"3c",X"2e",X"03",X"1a",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"9e",X"aa",X"98",X"0b",X"0b",X"0b",X"03",X"1a",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"2e",X"2f",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"62",X"51",X"18",X"8e",X"8e",X"41",X"51",X"62",X"51",X"15",X"cf",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"ed",X"2e",X"19",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"0b",X"3c",X"0b",X"17",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"92",X"61",X"0b",X"0b",X"0b",X"2f",X"03",X"1a",X"03",X"03",X"75",X"03",X"cc",X"0b",X"54",X"f0",X"6d",X"f0",X"6d",X"aa",X"12",X"aa",X"aa",X"aa",X"aa",X"54",X"3c",X"0b",X"aa",X"d6",X"d6",X"d6",X"2e",X"2e",X"0c",X"aa",X"0b",X"42",X"ea",X"1b",X"0b",X"00",X"6f",X"af",X"eb",X"f3",X"4e",X"f3",X"f3",X"ae",X"f3",X"ae",X"ae",X"39",X"ae",X"0b",X"1b",X"98",X"ed",X"54",X"2f",X"54",X"f0",X"54",X"2f",X"54",X"2f",X"54",X"f0",X"54",X"2f",X"54",X"f0",X"54",X"f0",X"0b",X"0b",X"2e",X"2e",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"2e",X"1b",X"0b",X"00",X"0b",X"87",X"39",X"39",X"ae",X"39",X"ae",X"82",X"ae",X"f3",X"f3",X"22",X"48",X"f3",X"4e",X"8b",X"eb",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"00",X"2e",X"19",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"70",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"60",X"aa",X"7c",X"aa",X"84",X"0b",X"0b",X"1b",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"2e",X"ed",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"f5",X"51",X"62",X"62",X"51",X"51",X"c7",X"8e",X"51",X"51",X"62",X"62",X"62",X"62",X"15",X"51",X"62",X"62",X"15",X"62",X"62",X"cf",X"62",X"2f",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"75",X"03",X"1a",X"71",X"19",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"27",X"19",X"71",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"0b",X"0b",X"3c",X"33",X"f0",X"6d",X"3f",X"6d",
    X"9e",X"aa",X"aa",X"aa",X"98",X"1b",X"0b",X"1b",X"61",X"03",X"19",X"71",X"19",X"b2",X"03",X"03",X"2e",X"3c",X"f0",X"6d",X"f0",X"6d",X"aa",X"60",X"aa",X"9e",X"54",X"0b",X"3c",X"0b",X"0b",X"a7",X"89",X"d6",X"d6",X"d6",X"2e",X"2e",X"ec",X"0c",X"0b",X"fc",X"0b",X"0b",X"8b",X"af",X"8b",X"4e",X"8b",X"f3",X"22",X"82",X"f3",X"ae",X"82",X"ae",X"82",X"39",X"39",X"f3",X"0b",X"1b",X"0b",X"ed",X"54",X"ed",X"54",X"f0",X"54",X"2f",X"54",X"ed",X"54",X"2f",X"0b",X"1b",X"0b",X"3c",X"0b",X"3c",X"0b",X"3c",X"2e",X"2e",X"19",X"03",X"71",X"19",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"2e",X"2e",X"1b",X"0b",X"0b",X"0b",X"39",X"4a",X"ae",X"82",X"ae",X"ae",X"ae",X"f3",X"f3",X"f3",X"4e",X"8b",X"4e",X"af",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"2e",X"03",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"aa",X"9e",X"aa",X"98",X"83",X"1b",X"0b",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"e5",X"2f",X"62",X"62",X"62",X"cf",X"15",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"1d",X"51",X"15",X"51",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"ed",X"2e",X"03",X"19",X"03",X"03",X"71",X"19",X"03",X"b2",X"19",X"71",X"03",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"1a",X"03",X"03",X"0b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"60",X"12",X"2c",X"61",X"0b",X"0b",X"0b",X"2f",X"03",X"b2",X"19",X"03",X"03",X"03",X"1a",X"ec",X"0b",X"54",X"6d",X"3f",X"6d",X"f0",X"aa",X"54",X"1b",X"3c",X"1b",X"2e",X"2e",X"3c",X"5f",X"68",X"0c",X"f8",X"d6",X"09",X"2e",X"2e",X"2e",X"ec",X"0b",X"0b",X"3c",X"4e",X"8b",X"4e",X"8b",X"f3",X"eb",X"f3",X"f3",X"ae",X"f3",X"ae",X"70",X"d1",X"ae",X"39",X"fb",X"d1",X"f3",X"0b",X"1b",X"0b",X"3c",X"54",X"ed",X"54",X"1b",X"0b",X"0b",X"3c",X"0b",X"0b",X"8b",X"af",X"6f",X"0b",X"1b",X"0b",X"0b",X"3c",X"0b",X"2e",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"75",X"03",X"21",X"2e",X"3c",X"0b",X"3c",X"0b",X"39",X"ae",X"ae",X"70",X"f3",X"ae",X"f3",X"6f",X"f3",X"4e",X"8b",X"8b",X"3c",X"0b",X"3c",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"91",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"12",X"aa",X"7c",X"aa",X"33",X"0b",X"0b",X"0b",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"27",X"b2",X"03",X"19",X"71",X"19",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"2e",X"54",X"62",X"15",X"51",X"62",X"62",X"cf",X"15",X"f5",X"51",X"62",X"cf",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"cf",X"62",X"51",X"62",X"62",X"cf",X"15",X"62",X"62",X"15",X"62",X"15",X"f5",X"ed",X"2e",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"e4",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"aa",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"79",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"2e",X"1b",X"0b",X"f0",X"6d",X"f0",X"54",X"0b",X"3c",X"0b",X"2e",X"2e",X"2e",X"2f",X"0b",X"a7",X"0c",X"0c",X"0c",X"f8",X"d6",X"d6",X"2e",X"2e",X"2e",X"a7",X"3c",X"0b",X"8b",X"af",X"8b",X"4e",X"8b",X"46",X"f3",X"22",X"f3",X"ae",X"ae",X"ae",X"82",X"39",X"39",X"39",X"d1",X"d1",X"f3",X"0b",X"3c",X"0b",X"0b",X"00",X"0b",X"0b",X"ae",X"39",X"39",X"39",X"fb",X"82",X"ae",X"70",X"4e",X"0b",X"0b",X"00",X"0b",X"0b",X"3c",X"2e",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"71",X"2e",X"1b",X"0b",X"00",X"0b",X"0b",X"82",X"ae",X"ae",X"f3",X"f3",X"22",X"48",X"f3",X"4e",X"eb",X"8b",X"1b",X"3b",X"3b",X"ce",X"10",X"ce",X"1c",X"10",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"70",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"3b",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"9e",X"aa",X"98",X"0b",X"0b",X"1b",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"2e",X"ed",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"15",X"62",X"cf",X"62",X"15",X"62",X"51",X"62",X"15",X"62",X"62",X"62",X"51",X"62",X"62",X"cf",X"62",X"51",X"62",X"62",X"51",X"79",X"2e",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"71",X"19",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"0b",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"3f",
    X"9e",X"7c",X"aa",X"60",X"61",X"0b",X"1b",X"0b",X"2f",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"b2",X"2e",X"3c",X"54",X"2f",X"0b",X"3c",X"2f",X"2e",X"2e",X"2e",X"2f",X"f0",X"73",X"1b",X"f0",X"a7",X"89",X"0c",X"0c",X"f8",X"f8",X"d6",X"2e",X"2e",X"2e",X"3c",X"0b",X"65",X"8b",X"4e",X"eb",X"f3",X"8b",X"f3",X"f3",X"ae",X"f3",X"ae",X"70",X"d1",X"82",X"d1",X"39",X"d1",X"d1",X"d1",X"0b",X"1b",X"0b",X"3c",X"0b",X"1b",X"b8",X"ff",X"d1",X"d1",X"4a",X"39",X"ae",X"ae",X"82",X"f3",X"48",X"3c",X"0b",X"0b",X"00",X"0b",X"00",X"2e",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"19",X"71",X"19",X"03",X"21",X"2e",X"0b",X"3c",X"0b",X"0b",X"0b",X"f3",X"ae",X"f3",X"f3",X"f3",X"4e",X"8b",X"4e",X"8b",X"3b",X"3b",X"10",X"b9",X"b9",X"b9",X"6c",X"07",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",X"60",X"aa",X"7c",X"aa",X"74",X"0b",X"1b",X"0b",X"19",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"19",X"03",X"71",X"27",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"d8",X"19",X"ec",X"f0",X"62",X"62",X"62",X"15",X"62",X"62",X"51",X"cf",X"62",X"62",X"51",X"62",X"51",X"62",X"cf",X"62",X"62",X"62",X"51",X"cf",X"15",X"51",X"62",X"62",X"51",X"15",X"62",X"62",X"51",X"62",X"62",X"2f",X"2e",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"1a",X"1b",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"0b",X"0b",X"77",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"03",X"cc",X"1b",X"0b",X"3c",X"0b",X"2e",X"2e",X"2e",X"1b",X"3c",X"73",X"d6",X"d6",X"aa",X"54",X"a7",X"5f",X"68",X"a7",X"aa",X"0c",X"f8",X"f8",X"d6",X"2e",X"0b",X"0b",X"af",X"4e",X"8b",X"4e",X"8b",X"f3",X"22",X"82",X"f3",X"ae",X"82",X"ae",X"ae",X"39",X"39",X"fb",X"39",X"d1",X"d1",X"f3",X"0b",X"3c",X"0b",X"0b",X"3c",X"39",X"d1",X"39",X"d1",X"39",X"39",X"39",X"ae",X"ae",X"ae",X"ae",X"8b",X"1b",X"1b",X"0b",X"0b",X"0b",X"0b",X"30",X"03",X"1a",X"03",X"03",X"b2",X"27",X"03",X"03",X"1a",X"03",X"b2",X"19",X"b2",X"03",X"1a",X"03",X"75",X"03",X"19",X"ec",X"2e",X"1b",X"0b",X"00",X"0b",X"f3",X"f3",X"22",X"8b",X"f3",X"4e",X"8b",X"af",X"3b",X"10",X"b9",X"2a",X"2a",X"2a",X"2a",X"b9",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"aa",X"9e",X"aa",X"98",X"1b",X"0b",X"0b",X"d8",X"b2",X"03",X"19",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"2e",X"54",X"51",X"62",X"51",X"cf",X"62",X"15",X"62",X"62",X"51",X"15",X"62",X"62",X"15",X"f5",X"51",X"62",X"51",X"62",X"62",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"61",X"2e",X"03",X"75",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"19",X"b2",X"27",X"19",X"03",X"75",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"03",X"19",X"7d",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"12",X"98",X"1b",X"0b",X"0b",X"2f",X"03",X"19",X"71",X"03",X"03",X"19",X"71",X"1a",X"03",X"cc",X"0b",X"21",X"2e",X"03",X"21",X"1b",X"54",X"6d",X"1b",X"d6",X"d6",X"e9",X"00",X"aa",X"a7",X"36",X"54",X"1b",X"3c",X"0c",X"0c",X"d6",X"0b",X"3c",X"1b",X"8b",X"8b",X"af",X"8b",X"f3",X"4e",X"f3",X"f3",X"ae",X"f3",X"ae",X"82",X"39",X"ae",X"39",X"39",X"d1",X"39",X"ff",X"d1",X"f3",X"0b",X"1b",X"0b",X"f3",X"d1",X"57",X"d1",X"39",X"d1",X"4a",X"39",X"39",X"ae",X"82",X"f3",X"f3",X"8b",X"0b",X"1b",X"1b",X"0b",X"3c",X"0b",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"71",X"19",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"ec",X"1b",X"0b",X"00",X"0b",X"0b",X"f3",X"f3",X"6f",X"af",X"8b",X"8b",X"cd",X"c1",X"2a",X"e3",X"e3",X"e3",X"2a",X"b9",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"12",X"aa",X"7c",X"aa",X"98",X"0b",X"0b",X"0b",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"19",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"19",X"2e",X"2f",X"62",X"62",X"15",X"62",X"51",X"f5",X"51",X"62",X"62",X"62",X"cf",X"62",X"51",X"62",X"15",X"62",X"15",X"62",X"51",X"62",X"51",X"62",X"cf",X"62",X"62",X"15",X"cf",X"15",X"62",X"62",X"62",X"2f",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"71",X"19",X"b2",X"27",X"19",X"03",X"03",X"b2",X"03",X"19",X"71",X"27",X"1a",X"03",X"19",X"b2",X"19",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"b2",X"83",X"3c",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"9e",X"aa",X"98",X"0b",X"1b",X"83",X"2f",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"03",X"19",X"03",X"30",X"19",X"03",X"2e",X"0b",X"54",X"aa",X"aa",X"6d",X"ed",X"73",X"4d",X"fc",X"6d",X"9e",X"a7",X"54",X"0b",X"73",X"1b",X"0c",X"54",X"fc",X"0b",X"0b",X"eb",X"4e",X"8b",X"4e",X"af",X"f3",X"22",X"f3",X"f3",X"ae",X"ae",X"ae",X"82",X"d1",X"39",X"4a",X"39",X"d1",X"d1",X"57",X"d1",X"0b",X"3c",X"0b",X"d1",X"57",X"d1",X"d1",X"d1",X"39",X"39",X"fb",X"ae",X"39",X"ae",X"ae",X"f3",X"f3",X"4e",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"2e",X"19",X"03",X"19",X"71",X"19",X"03",X"03",X"19",X"71",X"19",X"b2",X"27",X"03",X"1a",X"03",X"03",X"75",X"03",X"03",X"1a",X"2e",X"2e",X"1b",X"0b",X"3c",X"0b",X"00",X"3c",X"8b",X"4e",X"65",X"3b",X"bb",X"2a",X"2e",X"2e",X"e3",X"2a",X"b9",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"91",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"79",X"6d",X"f0",X"3f",X"6d",X"aa",X"aa",X"60",X"61",X"0b",X"0b",X"3c",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"d8",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"2e",X"ed",X"62",X"51",X"62",X"51",X"62",X"15",X"62",X"f5",X"51",X"62",X"51",X"15",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"51",X"54",X"2e",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"1b",X"0b",X"0b",X"53",X"6d",X"3f",X"6d",X"3f",
    X"aa",X"7c",X"aa",X"60",X"98",X"0b",X"1b",X"0b",X"79",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"b2",X"03",X"2e",X"3c",X"54",X"3f",X"aa",X"60",X"aa",X"6d",X"3c",X"0b",X"ea",X"1b",X"aa",X"9e",X"aa",X"54",X"f0",X"42",X"aa",X"42",X"d6",X"3c",X"0b",X"af",X"8b",X"eb",X"8b",X"f3",X"8b",X"f3",X"f3",X"ae",X"f3",X"ae",X"70",X"d1",X"82",X"39",X"d1",X"39",X"4a",X"57",X"d1",X"d1",X"57",X"0b",X"1b",X"d1",X"d1",X"d1",X"d1",X"39",X"fb",X"39",X"39",X"39",X"ae",X"ae",X"ae",X"ae",X"f3",X"f3",X"4e",X"0b",X"1b",X"0b",X"00",X"0b",X"0b",X"ec",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"75",X"03",X"03",X"b2",X"27",X"19",X"58",X"3b",X"3b",X"3b",X"3b",X"3b",X"33",X"3b",X"3b",X"2e",X"1b",X"0b",X"0b",X"0b",X"0b",X"3c",X"8b",X"3b",X"10",X"2a",X"2e",X"2e",X"e3",X"2a",X"b9",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"6d",X"aa",X"aa",X"60",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"03",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"2e",X"2f",X"62",X"62",X"62",X"62",X"51",X"62",X"51",X"15",X"62",X"62",X"62",X"62",X"cf",X"15",X"f5",X"51",X"cf",X"62",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"51",X"62",X"51",X"15",X"62",X"62",X"ed",X"2e",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"27",X"75",X"03",X"1a",X"03",X"19",X"03",X"75",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"0b",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"2f",X"03",X"b2",X"03",X"b2",X"27",X"03",X"1a",X"03",X"1a",X"03",X"03",X"2e",X"0b",X"2f",X"6d",X"f0",X"6d",X"aa",X"aa",X"aa",X"6d",X"ed",X"1b",X"0b",X"54",X"aa",X"7c",X"aa",X"0b",X"fc",X"ea",X"d6",X"2e",X"1b",X"0b",X"eb",X"48",X"4e",X"8b",X"4e",X"f3",X"22",X"82",X"f3",X"ae",X"ae",X"ae",X"82",X"39",X"ae",X"39",X"39",X"8a",X"39",X"d1",X"ff",X"d1",X"f3",X"0b",X"57",X"d1",X"ff",X"39",X"d1",X"39",X"d1",X"39",X"ae",X"39",X"82",X"70",X"f3",X"ae",X"f3",X"22",X"0b",X"3c",X"0b",X"0b",X"0b",X"3c",X"0b",X"2e",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"ad",X"3b",X"3b",X"3b",X"1c",X"10",X"ce",X"4e",X"eb",X"4e",X"3b",X"3b",X"3b",X"2e",X"1b",X"0b",X"3c",X"0b",X"1b",X"3b",X"1c",X"bb",X"b9",X"6c",X"2a",X"b9",X"07",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"70",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"92",X"aa",X"42",X"98",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"b2",X"27",X"19",X"71",X"27",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"2e",X"ed",X"62",X"51",X"62",X"15",X"cf",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"62",X"15",X"cf",X"62",X"15",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"cf",X"62",X"2f",X"2e",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"75",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"0b",X"0b",X"0b",X"3b",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"0d",X"60",X"61",X"0b",X"0b",X"0b",X"79",X"03",X"75",X"03",X"19",X"03",X"b2",X"19",X"71",X"19",X"03",X"75",X"2e",X"2f",X"0b",X"6d",X"f0",X"3f",X"6d",X"aa",X"9e",X"7c",X"f0",X"54",X"54",X"f0",X"aa",X"9e",X"aa",X"54",X"6d",X"d6",X"2e",X"3c",X"0b",X"0b",X"4e",X"eb",X"8b",X"af",X"f3",X"4e",X"f3",X"f3",X"ae",X"f3",X"ae",X"82",X"ae",X"ae",X"39",X"d1",X"4a",X"39",X"d1",X"d1",X"57",X"d1",X"d1",X"f3",X"d1",X"d1",X"57",X"d1",X"d1",X"87",X"39",X"4a",X"39",X"ae",X"ae",X"ae",X"82",X"82",X"f3",X"f3",X"f3",X"0b",X"1b",X"0b",X"3c",X"0b",X"0b",X"3c",X"2e",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1b",X"3b",X"10",X"1b",X"bb",X"3b",X"1c",X"10",X"1c",X"10",X"eb",X"8b",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"1c",X"bb",X"bb",X"bb",X"c1",X"bb",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"9e",X"aa",X"aa",X"6d",X"61",X"1b",X"0b",X"0b",X"03",X"b2",X"03",X"b2",X"d8",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"b2",X"19",X"03",X"03",X"1a",X"03",X"03",X"19",X"b2",X"2e",X"2f",X"62",X"62",X"51",X"62",X"62",X"15",X"cf",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"62",X"cf",X"15",X"62",X"51",X"62",X"51",X"62",X"51",X"77",X"2e",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"19",X"03",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"71",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"0b",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"7c",X"aa",X"98",X"0b",X"1b",X"0b",X"2f",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"21",X"54",X"2f",X"6d",X"6d",X"f0",X"6d",X"aa",X"9e",X"aa",X"7c",X"f0",X"aa",X"7c",X"aa",X"9e",X"f0",X"0b",X"2e",X"d6",X"fc",X"0b",X"3c",X"8b",X"4e",X"8b",X"4e",X"eb",X"f3",X"f3",X"f3",X"22",X"8b",X"00",X"1b",X"0b",X"65",X"ae",X"39",X"39",X"d1",X"39",X"ff",X"d1",X"d1",X"57",X"ae",X"d1",X"57",X"d1",X"39",X"d1",X"39",X"d1",X"39",X"ae",X"39",X"ae",X"70",X"ae",X"82",X"f3",X"f3",X"46",X"f3",X"0b",X"3c",X"0b",X"0b",X"3c",X"0b",X"0b",X"ec",X"03",X"19",X"03",X"03",X"1a",X"03",X"3b",X"3b",X"1c",X"bb",X"3b",X"e3",X"bb",X"3b",X"c1",X"10",X"ce",X"10",X"4e",X"eb",X"b6",X"74",X"b6",X"93",X"74",X"4e",X"8b",X"af",X"3b",X"3b",X"10",X"ce",X"1c",X"10",X"10",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"53",X"6d",X"79",X"6d",X"f0",X"aa",X"7c",X"aa",X"12",X"54",X"0b",X"0b",X"1b",X"03",X"19",X"03",X"19",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"03",X"19",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"2e",X"54",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"cf",X"62",X"51",X"62",X"62",X"62",X"51",X"15",X"62",X"62",X"cf",X"15",X"f5",X"62",X"62",X"62",X"ed",X"2e",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"27",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"71",X"03",X"1a",X"03",X"19",X"1b",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",
    X"aa",X"9e",X"aa",X"9e",X"98",X"0b",X"0b",X"1b",X"61",X"03",X"19",X"03",X"75",X"03",X"03",X"03",X"1a",X"03",X"03",X"03",X"19",X"03",X"21",X"1b",X"54",X"f0",X"6d",X"3f",X"6d",X"f0",X"9e",X"aa",X"60",X"aa",X"12",X"aa",X"7c",X"f0",X"0b",X"d6",X"0b",X"2e",X"3c",X"0b",X"65",X"8b",X"af",X"8b",X"f3",X"4e",X"f3",X"22",X"f3",X"1b",X"0b",X"0b",X"00",X"0b",X"0b",X"4a",X"39",X"d1",X"d1",X"d1",X"d1",X"57",X"d1",X"57",X"d1",X"d1",X"57",X"d1",X"d1",X"39",X"4a",X"39",X"4a",X"ae",X"82",X"ae",X"ae",X"f3",X"ae",X"f3",X"f3",X"f3",X"4e",X"0b",X"1b",X"0b",X"3c",X"0b",X"3c",X"2e",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"10",X"bb",X"07",X"3b",X"e3",X"2e",X"bb",X"3b",X"3b",X"c1",X"10",X"1c",X"4e",X"8b",X"9a",X"c7",X"c7",X"c7",X"4c",X"74",X"3b",X"4e",X"eb",X"3b",X"3b",X"3b",X"3b",X"3b",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"70",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"91",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"60",X"aa",X"9e",X"aa",X"74",X"0b",X"1b",X"0b",X"19",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"d8",X"19",X"71",X"19",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"e5",X"2f",X"62",X"62",X"15",X"cf",X"62",X"62",X"51",X"62",X"cf",X"15",X"62",X"cf",X"15",X"62",X"62",X"15",X"62",X"62",X"15",X"62",X"cf",X"62",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"98",X"2e",X"03",X"b2",X"03",X"19",X"03",X"75",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"ad",X"1b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"aa",X"33",X"1b",X"0b",X"0b",X"2f",X"03",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"2e",X"3c",X"54",X"f0",X"6d",X"f0",X"6d",X"f0",X"6d",X"aa",X"9e",X"aa",X"6d",X"f0",X"6d",X"2f",X"0b",X"ec",X"2e",X"0b",X"1b",X"8b",X"4e",X"8b",X"4e",X"8b",X"f3",X"f3",X"f3",X"82",X"0b",X"0b",X"3c",X"0b",X"1b",X"1b",X"0b",X"39",X"d1",X"39",X"d1",X"ff",X"d1",X"d1",X"d1",X"57",X"d1",X"d1",X"39",X"1f",X"39",X"d1",X"39",X"ae",X"39",X"ae",X"ae",X"82",X"ae",X"f3",X"f3",X"22",X"f3",X"f3",X"6f",X"3c",X"0b",X"0b",X"0b",X"0b",X"3c",X"2e",X"7f",X"e3",X"e3",X"6c",X"1c",X"3b",X"3b",X"3b",X"bb",X"3b",X"e3",X"2e",X"2e",X"bb",X"10",X"3b",X"c1",X"10",X"22",X"af",X"4c",X"2e",X"2e",X"2e",X"af",X"8b",X"23",X"3b",X"46",X"8b",X"3b",X"03",X"3b",X"74",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"aa",X"7c",X"aa",X"98",X"1b",X"0b",X"0b",X"03",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"27",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"2e",X"2f",X"f5",X"51",X"62",X"62",X"15",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"51",X"62",X"15",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"15",X"2f",X"2e",X"03",X"75",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"75",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"9e",X"7c",X"61",X"0b",X"0b",X"1b",X"61",X"03",X"75",X"03",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"2e",X"3c",X"0b",X"2f",X"6d",X"6d",X"f0",X"3f",X"6d",X"f0",X"6d",X"3f",X"6d",X"2f",X"0b",X"2e",X"1a",X"03",X"cc",X"3c",X"0b",X"af",X"4e",X"8b",X"f3",X"4e",X"f3",X"f3",X"22",X"0b",X"0b",X"3c",X"0b",X"b2",X"03",X"0b",X"3c",X"4a",X"57",X"d1",X"57",X"d1",X"57",X"57",X"d1",X"d1",X"ff",X"d1",X"39",X"39",X"4a",X"39",X"39",X"ae",X"ae",X"70",X"ae",X"f3",X"ae",X"f3",X"f3",X"f3",X"6f",X"af",X"0b",X"1b",X"0b",X"00",X"3c",X"0b",X"0b",X"2e",X"3b",X"e3",X"2e",X"2e",X"e3",X"6c",X"1c",X"3b",X"3b",X"e3",X"2e",X"2e",X"2e",X"e3",X"bb",X"3b",X"bb",X"10",X"22",X"8b",X"23",X"c7",X"6f",X"3b",X"3b",X"8b",X"74",X"17",X"d7",X"3b",X"3b",X"3b",X"3b",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"60",X"aa",X"9e",X"54",X"0b",X"0b",X"1b",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"75",X"03",X"2e",X"f0",X"15",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"15",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"51",X"62",X"15",X"cf",X"62",X"f0",X"2e",X"b2",X"03",X"03",X"19",X"03",X"03",X"75",X"03",X"19",X"71",X"19",X"03",X"b2",X"19",X"71",X"27",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"d8",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"03",X"0b",X"0b",X"0b",X"17",X"f0",X"6d",X"3f",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"2f",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"19",X"03",X"19",X"b2",X"2e",X"1b",X"0b",X"2f",X"6d",X"f0",X"6d",X"6d",X"f0",X"6d",X"f0",X"54",X"1b",X"0b",X"cc",X"03",X"03",X"2e",X"0b",X"0b",X"65",X"8b",X"af",X"8b",X"22",X"f3",X"22",X"f3",X"1b",X"3c",X"0b",X"0b",X"03",X"19",X"71",X"1b",X"0b",X"39",X"d1",X"d1",X"d1",X"d1",X"d1",X"d1",X"57",X"d1",X"39",X"d1",X"d1",X"39",X"d1",X"82",X"39",X"ae",X"ae",X"ae",X"b7",X"b8",X"f3",X"46",X"f3",X"f3",X"4e",X"8b",X"3c",X"0b",X"0b",X"0b",X"0b",X"3c",X"0b",X"2e",X"3b",X"e3",X"2e",X"2e",X"2e",X"2e",X"e3",X"e3",X"e3",X"2e",X"2e",X"2e",X"2e",X"2e",X"e3",X"3b",X"1c",X"46",X"eb",X"3b",X"b6",X"af",X"2e",X"3b",X"4e",X"74",X"3b",X"46",X"8b",X"3b",X"3b",X"ce",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"3b",X"f0",X"6d",X"f0",X"6d",X"12",X"aa",X"7c",X"aa",X"84",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"03",X"19",X"03",X"75",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"2e",X"1a",X"62",X"51",X"62",X"62",X"15",X"cf",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"cf",X"15",X"51",X"cf",X"62",X"15",X"51",X"62",X"62",X"cf",X"15",X"62",X"cf",X"62",X"62",X"62",X"51",X"62",X"28",X"2e",X"03",X"19",X"b2",X"19",X"71",X"19",X"71",X"03",X"b2",X"19",X"03",X"75",X"03",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"03",X"b2",X"03",X"b2",X"19",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"79",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"cc",X"2e",X"1b",X"0b",X"2f",X"6d",X"f0",X"6d",X"f0",X"54",X"1b",X"0b",X"ec",X"03",X"03",X"1a",X"ec",X"0b",X"1b",X"8b",X"4e",X"8b",X"af",X"8b",X"f3",X"f3",X"f3",X"8b",X"1b",X"0b",X"00",X"19",X"71",X"19",X"3c",X"0b",X"d1",X"d1",X"57",X"d1",X"57",X"d1",X"57",X"d1",X"d1",X"ff",X"39",X"4a",X"39",X"39",X"fb",X"82",X"ae",X"70",X"ae",X"82",X"70",X"f3",X"f3",X"f3",X"6f",X"f3",X"4e",X"8b",X"00",X"0b",X"00",X"0b",X"3c",X"0b",X"ec",X"3b",X"3b",X"e3",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"e3",X"3b",X"d7",X"8b",X"3b",X"3b",X"ef",X"8b",X"af",X"74",X"3b",X"33",X"eb",X"22",X"3b",X"10",X"1c",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"aa",X"9e",X"aa",X"98",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"03",X"19",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"ec",X"1a",X"15",X"f5",X"51",X"62",X"62",X"51",X"f5",X"62",X"15",X"cf",X"62",X"51",X"62",X"51",X"62",X"62",X"15",X"62",X"cf",X"62",X"62",X"15",X"51",X"62",X"62",X"15",X"f5",X"51",X"62",X"62",X"62",X"75",X"2e",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"19",X"b2",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"27",X"19",X"03",X"19",X"03",X"0b",X"0b",X"1b",X"33",X"f0",X"6d",X"f0",X"3f",
    X"aa",X"7c",X"aa",X"aa",X"84",X"0b",X"0b",X"0b",X"2f",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"21",X"2e",X"1b",X"0b",X"3c",X"1b",X"3c",X"0b",X"30",X"cc",X"1a",X"03",X"1a",X"03",X"e5",X"3c",X"0b",X"65",X"8b",X"4e",X"8b",X"f3",X"4e",X"f3",X"f3",X"22",X"0b",X"0b",X"3c",X"0b",X"03",X"1a",X"03",X"0b",X"0b",X"d1",X"57",X"d1",X"d1",X"57",X"d1",X"d1",X"57",X"d1",X"d1",X"39",X"4a",X"39",X"ae",X"39",X"ae",X"82",X"ae",X"ae",X"f3",X"ae",X"f3",X"22",X"f3",X"48",X"f3",X"6f",X"1b",X"0b",X"0b",X"00",X"0b",X"0b",X"0b",X"3b",X"c1",X"3b",X"b9",X"e3",X"2e",X"2e",X"2e",X"2e",X"2e",X"e3",X"e3",X"e3",X"2e",X"2e",X"2e",X"e3",X"3b",X"4e",X"3b",X"3b",X"3b",X"3b",X"33",X"3b",X"3b",X"3b",X"3b",X"46",X"3b",X"1c",X"bb",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"33",X"79",X"6d",X"6d",X"f0",X"60",X"aa",X"7c",X"9e",X"98",X"0b",X"1b",X"0b",X"03",X"b2",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"27",X"75",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"cc",X"03",X"1a",X"15",X"62",X"51",X"62",X"62",X"15",X"51",X"62",X"62",X"15",X"62",X"62",X"62",X"62",X"51",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"15",X"62",X"51",X"15",X"1a",X"ec",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"0b",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"6d",
    X"9e",X"aa",X"7c",X"9e",X"98",X"0b",X"83",X"1b",X"2f",X"19",X"03",X"b2",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"75",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"ec",X"2e",X"2e",X"2e",X"2e",X"2e",X"03",X"03",X"03",X"03",X"03",X"b2",X"03",X"2e",X"1b",X"0b",X"4e",X"8b",X"4e",X"6f",X"f3",X"f3",X"46",X"f3",X"0b",X"3c",X"0b",X"0b",X"0b",X"3c",X"03",X"0b",X"00",X"d1",X"d1",X"57",X"d1",X"d1",X"d1",X"57",X"d1",X"39",X"1b",X"0b",X"3c",X"0b",X"39",X"82",X"ae",X"ae",X"70",X"ae",X"ae",X"f3",X"f3",X"82",X"f3",X"22",X"af",X"8b",X"af",X"0b",X"1b",X"0b",X"0b",X"00",X"3b",X"3b",X"bb",X"07",X"3b",X"3b",X"e3",X"2e",X"2e",X"2e",X"2e",X"e3",X"3b",X"3b",X"b9",X"e3",X"2e",X"2e",X"e3",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"22",X"3b",X"c1",X"07",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"70",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"3f",X"f0",X"6d",X"aa",X"60",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"03",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"75",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"2e",X"19",X"1a",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"15",X"62",X"51",X"62",X"51",X"62",X"62",X"51",X"62",X"51",X"51",X"62",X"62",X"62",X"51",X"62",X"75",X"19",X"2e",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"27",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"71",X"19",X"03",X"03",X"1a",X"1b",X"0b",X"0b",X"98",X"f0",X"6d",X"f0",X"3f",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"79",X"03",X"b2",X"19",X"03",X"75",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"b2",X"19",X"b2",X"19",X"03",X"19",X"2e",X"00",X"0b",X"af",X"8b",X"af",X"f3",X"6f",X"f3",X"f3",X"f3",X"f3",X"f3",X"1b",X"0b",X"00",X"0b",X"0b",X"1b",X"0b",X"0b",X"d1",X"d1",X"57",X"d1",X"57",X"d1",X"d1",X"1b",X"0b",X"0b",X"3c",X"0b",X"3c",X"0b",X"ae",X"82",X"ae",X"ae",X"f3",X"ae",X"f3",X"22",X"f3",X"8b",X"f3",X"8b",X"4e",X"0b",X"00",X"0b",X"1b",X"0b",X"3b",X"10",X"c1",X"b9",X"b9",X"10",X"ad",X"6c",X"2e",X"2e",X"2e",X"e3",X"3b",X"2a",X"3b",X"3b",X"b9",X"e3",X"e3",X"e3",X"3b",X"3b",X"3b",X"74",X"74",X"3b",X"3b",X"3b",X"3b",X"46",X"3b",X"bb",X"b9",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"f4",X"91",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"aa",X"aa",X"9e",X"98",X"1b",X"0b",X"0b",X"19",X"71",X"19",X"b2",X"27",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"d8",X"19",X"03",X"19",X"b2",X"19",X"71",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"2e",X"03",X"1a",X"75",X"62",X"62",X"15",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"51",X"62",X"62",X"62",X"51",X"62",X"62",X"62",X"62",X"62",X"62",X"15",X"51",X"75",X"03",X"b2",X"2e",X"03",X"b2",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"b2",X"19",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"03",X"19",X"03",X"b2",X"27",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"0b",X"0b",X"0b",X"3b",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"9e",X"98",X"0b",X"1b",X"0b",X"2f",X"19",X"03",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"b2",X"2e",X"1b",X"0b",X"8b",X"af",X"6f",X"8b",X"f3",X"22",X"f3",X"f3",X"ae",X"f3",X"82",X"48",X"0b",X"3c",X"0b",X"00",X"0b",X"1b",X"39",X"1f",X"57",X"d1",X"d1",X"57",X"d1",X"0b",X"0b",X"00",X"0b",X"0b",X"03",X"0b",X"0b",X"82",X"ae",X"70",X"ae",X"f3",X"f3",X"f3",X"82",X"22",X"4e",X"f3",X"6f",X"af",X"0b",X"0b",X"00",X"0b",X"3b",X"ce",X"6c",X"2a",X"2a",X"2a",X"2a",X"3b",X"b9",X"e3",X"2e",X"e3",X"3b",X"2a",X"2a",X"b9",X"3b",X"3b",X"3b",X"b9",X"e3",X"3b",X"74",X"af",X"4e",X"74",X"3b",X"3b",X"3b",X"22",X"53",X"b9",X"b9",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"f3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"7c",X"9e",X"7c",X"61",X"0b",X"0b",X"1b",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"75",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"71",X"19",X"03",X"b2",X"19",X"03",X"1a",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"e5",X"03",X"1a",X"03",X"f0",X"f0",X"f0",X"f0",X"f0",X"98",X"f0",X"f0",X"98",X"f0",X"f0",X"2f",X"f0",X"f0",X"98",X"f0",X"2f",X"f0",X"f0",X"f0",X"1a",X"19",X"03",X"1a",X"2e",X"03",X"b2",X"19",X"03",X"75",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"b2",X"cd",X"0b",X"1b",X"33",X"6d",X"3f",X"6d",X"f0",
    X"9e",X"aa",X"60",X"aa",X"98",X"0b",X"83",X"0b",X"79",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"03",X"b2",X"27",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"2e",X"00",X"0b",X"65",X"4e",X"af",X"f3",X"4e",X"f3",X"f3",X"22",X"f3",X"ae",X"ae",X"ae",X"82",X"8b",X"1b",X"0b",X"0b",X"00",X"0b",X"39",X"d1",X"d1",X"ff",X"d1",X"d1",X"0b",X"1b",X"0b",X"0b",X"03",X"03",X"b2",X"1b",X"0b",X"ae",X"ae",X"ae",X"ae",X"f3",X"f3",X"22",X"f3",X"f3",X"8b",X"af",X"6f",X"1b",X"0b",X"3c",X"0b",X"3b",X"c1",X"2a",X"2a",X"e3",X"e3",X"e3",X"e3",X"3b",X"3b",X"6c",X"e3",X"3b",X"2a",X"2a",X"b9",X"bb",X"1c",X"46",X"3b",X"3b",X"74",X"8b",X"3b",X"3b",X"4e",X"74",X"3b",X"8b",X"d7",X"3b",X"b9",X"2a",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"70",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"4a",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"9e",X"aa",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"b2",X"19",X"03",X"75",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"cc",X"2e",X"2e",X"ec",X"2e",X"2e",X"2e",X"2e",X"ec",X"2e",X"2e",X"ec",X"2e",X"2e",X"2e",X"2e",X"ec",X"2e",X"2e",X"e5",X"2e",X"ec",X"2e",X"2e",X"30",X"2e",X"2e",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"2f",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"2e",X"1b",X"0b",X"8b",X"8b",X"af",X"f3",X"f3",X"46",X"f3",X"ae",X"f3",X"ae",X"70",X"d1",X"f3",X"fb",X"8b",X"1b",X"0b",X"0b",X"ff",X"d1",X"d1",X"57",X"d1",X"57",X"0b",X"3c",X"0b",X"3c",X"03",X"03",X"03",X"75",X"3c",X"82",X"ae",X"70",X"f3",X"ae",X"f3",X"f3",X"82",X"6f",X"f3",X"4e",X"8b",X"4e",X"0b",X"0b",X"0b",X"3b",X"bb",X"2a",X"e3",X"e3",X"e3",X"e3",X"e3",X"e3",X"1c",X"3b",X"b9",X"3b",X"2a",X"2a",X"b9",X"07",X"10",X"22",X"af",X"93",X"4c",X"4e",X"2e",X"3b",X"8b",X"74",X"3b",X"46",X"d7",X"3b",X"b9",X"2a",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"82",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"f3",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"9e",X"7c",X"aa",X"84",X"0b",X"0b",X"1b",X"03",X"19",X"71",X"03",X"19",X"b2",X"19",X"71",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"75",X"03",X"03",X"b2",X"19",X"b2",X"27",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"19",X"71",X"19",X"71",X"19",X"71",X"19",X"03",X"b2",X"03",X"75",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"9e",X"aa",X"60",X"61",X"0b",X"1b",X"0b",X"77",X"03",X"1a",X"03",X"75",X"03",X"71",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"19",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"75",X"03",X"75",X"03",X"cc",X"3c",X"0b",X"eb",X"4e",X"f3",X"4e",X"f3",X"f3",X"f3",X"f3",X"ae",X"ae",X"82",X"ae",X"39",X"39",X"4a",X"39",X"22",X"f3",X"39",X"d1",X"57",X"d1",X"d1",X"d1",X"0b",X"1b",X"0b",X"0b",X"03",X"03",X"b2",X"27",X"1b",X"0b",X"ae",X"82",X"ae",X"f3",X"f3",X"f3",X"22",X"f3",X"4e",X"8b",X"af",X"8b",X"3c",X"0b",X"00",X"3b",X"c1",X"2a",X"e3",X"e3",X"e3",X"e3",X"e3",X"e3",X"e3",X"e3",X"3b",X"17",X"2a",X"b9",X"bb",X"1c",X"22",X"8b",X"23",X"4c",X"c7",X"2e",X"8b",X"af",X"2e",X"b6",X"3b",X"22",X"8b",X"cd",X"2a",X"2a",X"00",X"00",X"f4",X"00",X"2e",X"f4",X"82",X"3c",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3c",X"70",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",X"7c",X"aa",X"9e",X"aa",X"98",X"0b",X"0b",X"1b",X"19",X"71",X"19",X"19",X"b2",X"03",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"71",X"19",X"71",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"b2",X"19",X"03",X"03",X"75",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"d8",X"03",X"19",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"71",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"75",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"0b",X"3c",X"0b",X"3b",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"0b",X"0b",X"79",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"19",X"03",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"cc",X"0b",X"1b",X"0b",X"65",X"8b",X"f3",X"f3",X"22",X"f3",X"ae",X"f3",X"ae",X"ae",X"39",X"ae",X"39",X"d1",X"87",X"39",X"39",X"8a",X"d1",X"d1",X"57",X"d1",X"57",X"f3",X"0b",X"3c",X"0b",X"00",X"0b",X"03",X"03",X"b2",X"1b",X"82",X"ae",X"f3",X"ae",X"f3",X"22",X"f3",X"48",X"f3",X"6f",X"af",X"6f",X"af",X"0b",X"0b",X"cd",X"bb",X"2a",X"e3",X"2e",X"2e",X"e3",X"e3",X"e3",X"e3",X"e3",X"2a",X"2a",X"2a",X"b9",X"ce",X"46",X"4e",X"74",X"4c",X"c7",X"c7",X"2e",X"2e",X"2e",X"c7",X"74",X"3b",X"46",X"1c",X"3b",X"2a",X"e3",X"00",X"00",X"fb",X"00",X"2e",X"fb",X"82",X"82",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"f3",X"82",X"fb",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"12",X"aa",X"aa",X"7c",X"61",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"71",X"03",X"03",X"19",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"27",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"03",X"03",X"19",X"03",X"b2",X"27",X"1a",X"03",X"03",X"1a",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"b2",X"19",X"b2",X"27",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"b2",X"d8",X"03",X"0b",X"0b",X"0b",X"98",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"9e",X"aa",X"98",X"0b",X"1b",X"0b",X"79",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"75",X"03",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"75",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"03",X"cc",X"3c",X"0b",X"0b",X"f3",X"4e",X"f3",X"f3",X"f3",X"f3",X"ae",X"ae",X"70",X"ae",X"39",X"39",X"4a",X"39",X"d1",X"d1",X"39",X"d1",X"57",X"d1",X"57",X"d1",X"ae",X"0b",X"0b",X"1b",X"0b",X"0b",X"00",X"0b",X"19",X"3c",X"0b",X"ae",X"ae",X"f3",X"f3",X"82",X"f3",X"22",X"af",X"f3",X"6f",X"af",X"6f",X"1b",X"0b",X"3b",X"9b",X"2a",X"2e",X"2e",X"2e",X"2e",X"e3",X"e3",X"e3",X"e3",X"2a",X"2a",X"b9",X"bb",X"22",X"8b",X"3b",X"74",X"4c",X"c7",X"2e",X"2e",X"2e",X"2e",X"4c",X"6a",X"22",X"8b",X"cd",X"3b",X"2a",X"2e",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"f4",X"82",X"70",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"70",X"f4",X"91",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"3f",X"6d",X"aa",X"12",X"aa",X"98",X"0b",X"0b",X"0b",X"19",X"03",X"75",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"03",X"19",X"b2",X"27",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"d8",X"75",X"03",X"71",X"19",X"b2",X"27",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"b2",X"19",X"03",X"71",X"19",X"71",X"19",X"03",X"71",X"19",X"b2",X"d8",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"19",X"0b",X"1b",X"0b",X"3b",X"f0",X"6d",X"3f",X"6d",
    X"aa",X"7c",X"aa",X"92",X"61",X"0b",X"0b",X"0b",X"2f",X"03",X"1a",X"03",X"03",X"03",X"b2",X"27",X"03",X"1a",X"03",X"75",X"03",X"19",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"1a",X"03",X"2e",X"1b",X"3c",X"0b",X"0b",X"f3",X"b8",X"f3",X"ae",X"82",X"82",X"ae",X"39",X"ae",X"39",X"d1",X"39",X"39",X"4a",X"d1",X"57",X"d1",X"d1",X"d1",X"d1",X"57",X"39",X"ae",X"f3",X"0b",X"1b",X"0b",X"3c",X"0b",X"0b",X"00",X"82",X"f3",X"ae",X"f3",X"22",X"f3",X"8b",X"f3",X"4e",X"8b",X"af",X"8b",X"af",X"0b",X"3b",X"10",X"2a",X"2e",X"2e",X"2e",X"2e",X"e3",X"e3",X"e3",X"2a",X"2a",X"b9",X"bb",X"d7",X"af",X"3b",X"74",X"4c",X"c7",X"9a",X"2e",X"2e",X"2e",X"4c",X"74",X"3b",X"d7",X"4e",X"17",X"9f",X"2e",X"2e",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"fb",X"f4",X"91",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"91",X"f4",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"6d",X"aa",X"aa",X"2c",X"aa",X"84",X"0b",X"1b",X"0b",X"03",X"b2",X"27",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"27",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"75",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"0b",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"1b",X"1b",X"61",X"03",X"19",X"71",X"19",X"b2",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"b2",X"27",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"2e",X"2e",X"1b",X"3c",X"0b",X"00",X"f3",X"f3",X"ae",X"ae",X"ae",X"ae",X"39",X"4a",X"39",X"39",X"4a",X"57",X"39",X"d1",X"d1",X"57",X"d1",X"57",X"d1",X"d1",X"57",X"d1",X"ae",X"f3",X"0b",X"1b",X"0b",X"3c",X"0b",X"0b",X"ae",X"f3",X"f3",X"f3",X"82",X"22",X"8b",X"f3",X"4e",X"8b",X"4e",X"8b",X"3c",X"3b",X"10",X"b9",X"2a",X"2e",X"2e",X"e3",X"e3",X"e3",X"e3",X"2a",X"b9",X"97",X"d7",X"8b",X"3b",X"3b",X"ef",X"4c",X"9a",X"c7",X"c7",X"4c",X"74",X"74",X"3b",X"d7",X"af",X"10",X"3b",X"bb",X"2e",X"2e",X"00",X"00",X"f4",X"00",X"2e",X"fb",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"91",X"f4",X"fb",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"4f",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"12",X"aa",X"12",X"aa",X"98",X"0b",X"0b",X"0b",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"03",X"1a",X"03",X"71",X"75",X"03",X"1a",X"03",X"71",X"19",X"03",X"19",X"03",X"19",X"03",X"b2",X"27",X"1a",X"03",X"19",X"b2",X"03",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"06",X"19",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"b2",X"03",X"1a",X"03",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"7c",X"9e",X"6d",X"ba",X"0b",X"0b",X"0b",X"2f",X"03",X"b2",X"19",X"03",X"03",X"03",X"19",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"19",X"b2",X"27",X"19",X"b2",X"27",X"19",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"2e",X"2e",X"1b",X"0b",X"0b",X"00",X"f3",X"82",X"ae",X"39",X"ae",X"39",X"d1",X"4a",X"39",X"39",X"1f",X"57",X"d1",X"d1",X"57",X"d1",X"d1",X"57",X"d1",X"d1",X"d1",X"39",X"f3",X"0b",X"0b",X"1b",X"0b",X"3c",X"82",X"ae",X"f3",X"f3",X"22",X"f3",X"f3",X"6f",X"af",X"8b",X"eb",X"8b",X"3c",X"ad",X"3b",X"bb",X"2a",X"6b",X"e3",X"e3",X"e3",X"e3",X"2a",X"2a",X"b9",X"d7",X"af",X"af",X"3b",X"3b",X"3b",X"ef",X"6a",X"74",X"74",X"74",X"3b",X"3b",X"46",X"22",X"8b",X"3b",X"3b",X"bb",X"b9",X"2e",X"00",X"00",X"fb",X"00",X"2e",X"f4",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"2c",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"19",X"03",X"1a",X"03",X"03",X"19",X"03",X"1a",X"03",X"03",X"75",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"19",X"03",X"b2",X"d8",X"03",X"19",X"71",X"75",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"75",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"03",X"03",X"03",X"03",X"b2",X"03",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"83",X"3c",X"0b",X"53",X"6d",X"f0",X"6d",X"3f",
    X"9e",X"aa",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"79",X"03",X"19",X"03",X"b2",X"19",X"b2",X"27",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"03",X"1a",X"ec",X"2e",X"1b",X"0b",X"0b",X"00",X"f3",X"82",X"39",X"4a",X"39",X"39",X"d1",X"d1",X"39",X"d1",X"d1",X"57",X"d1",X"d1",X"57",X"d1",X"d1",X"d1",X"39",X"4a",X"39",X"ae",X"f3",X"0b",X"0b",X"1b",X"8b",X"f3",X"ae",X"f3",X"f3",X"46",X"8b",X"f3",X"4e",X"8b",X"4e",X"8b",X"af",X"1b",X"3b",X"1c",X"6c",X"2a",X"e3",X"6b",X"e3",X"e3",X"2a",X"b9",X"af",X"d7",X"8b",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"d7",X"d7",X"8b",X"ce",X"3b",X"1c",X"10",X"c1",X"6c",X"00",X"00",X"f4",X"3c",X"8f",X"4f",X"fb",X"91",X"00",X"3c",X"3c",X"00",X"fb",X"f4",X"fb",X"91",X"00",X"3c",X"3c",X"fb",X"f4",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5d",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"12",X"aa",X"92",X"61",X"0b",X"0b",X"0b",X"03",X"b2",X"03",X"19",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"03",X"19",X"03",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"19",X"71",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"19",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"92",X"61",X"0b",X"0b",X"0b",X"2f",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"cc",X"e5",X"1b",X"0b",X"00",X"0b",X"f3",X"39",X"d1",X"4a",X"39",X"d1",X"d1",X"d1",X"57",X"d1",X"d1",X"57",X"d1",X"d1",X"57",X"39",X"8a",X"39",X"fb",X"39",X"ae",X"39",X"ae",X"0b",X"0b",X"82",X"f3",X"ae",X"f3",X"f3",X"f3",X"4e",X"8b",X"af",X"8b",X"4e",X"8b",X"0b",X"3b",X"10",X"c1",X"2a",X"e3",X"e3",X"e3",X"2a",X"2a",X"b9",X"4e",X"f3",X"4e",X"17",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"33",X"17",X"46",X"d7",X"eb",X"10",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"f4",X"3c",X"a4",X"8f",X"a4",X"3c",X"f4",X"4f",X"f4",X"fb",X"a4",X"8f",X"8f",X"3c",X"91",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"3b",X"f0",X"6d",X"3f",X"6d",X"aa",X"2c",X"aa",X"aa",X"ba",X"0b",X"0b",X"1b",X"03",X"1a",X"03",X"b2",X"03",X"03",X"75",X"03",X"03",X"03",X"1a",X"03",X"03",X"1a",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"03",X"75",X"03",X"b2",X"19",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"03",X"b2",X"27",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"83",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"9e",X"aa",X"98",X"0b",X"0b",X"1b",X"61",X"03",X"75",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"75",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"cc",X"2e",X"0b",X"3c",X"0b",X"00",X"82",X"39",X"39",X"d1",X"39",X"ff",X"d1",X"d1",X"57",X"d1",X"57",X"d1",X"d1",X"d1",X"39",X"39",X"39",X"39",X"39",X"ae",X"ae",X"ae",X"ae",X"ae",X"ae",X"f3",X"f3",X"82",X"6f",X"f3",X"8b",X"4e",X"eb",X"8b",X"af",X"0b",X"3b",X"3b",X"c1",X"9f",X"2a",X"2a",X"2a",X"2a",X"2a",X"b9",X"af",X"d7",X"46",X"8b",X"53",X"3b",X"3b",X"3b",X"17",X"3b",X"22",X"46",X"22",X"8b",X"10",X"3b",X"3b",X"3b",X"4c",X"4c",X"4c",X"3b",X"00",X"00",X"f4",X"3c",X"8f",X"4f",X"fb",X"a4",X"8f",X"a4",X"8f",X"3c",X"fb",X"f4",X"f4",X"fb",X"8f",X"a4",X"a4",X"a4",X"3c",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"12",X"aa",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"19",X"03",X"1a",X"03",X"03",X"1a",X"71",X"19",X"71",X"1a",X"03",X"71",X"19",X"03",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"b2",X"19",X"71",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"71",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"d8",X"75",X"03",X"71",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"3c",X"0b",X"0b",X"53",X"6d",X"3f",X"6d",X"f0",
    X"aa",X"aa",X"7c",X"aa",X"84",X"0b",X"0b",X"0b",X"2f",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"21",X"2e",X"1b",X"0b",X"0b",X"00",X"ae",X"39",X"d1",X"d1",X"ff",X"d1",X"d1",X"d1",X"ff",X"d1",X"57",X"d1",X"d1",X"d1",X"39",X"fb",X"ae",X"39",X"ae",X"70",X"ae",X"70",X"f3",X"ae",X"f3",X"22",X"f3",X"af",X"4e",X"8b",X"4e",X"8b",X"cd",X"3b",X"3b",X"3b",X"10",X"bb",X"b9",X"fa",X"2a",X"2a",X"b9",X"9f",X"b9",X"af",X"d7",X"d7",X"22",X"22",X"46",X"22",X"46",X"22",X"46",X"eb",X"4e",X"1c",X"3b",X"3b",X"3b",X"4c",X"9a",X"c7",X"4c",X"4c",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"f4",X"8f",X"a4",X"8f",X"a4",X"3c",X"91",X"f4",X"4f",X"91",X"a4",X"8f",X"a4",X"8f",X"3c",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"60",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"19",X"03",X"75",X"03",X"b2",X"19",X"71",X"19",X"03",X"19",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"71",X"19",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"27",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"1a",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"19",X"b2",X"19",X"03",X"03",X"0b",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"60",X"aa",X"12",X"aa",X"98",X"0b",X"83",X"3c",X"2f",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"75",X"03",X"03",X"b2",X"03",X"75",X"03",X"19",X"b2",X"27",X"19",X"03",X"19",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"b2",X"27",X"19",X"03",X"2e",X"2e",X"1b",X"0b",X"0b",X"00",X"ae",X"39",X"d1",X"d1",X"57",X"d1",X"57",X"d1",X"d1",X"ff",X"39",X"1f",X"39",X"39",X"39",X"ae",X"ae",X"ae",X"ae",X"82",X"ae",X"f3",X"f3",X"f3",X"8b",X"22",X"8b",X"8b",X"af",X"3b",X"3b",X"4e",X"af",X"6f",X"3b",X"1c",X"bb",X"b9",X"b9",X"bb",X"9f",X"b9",X"b9",X"bb",X"4e",X"8b",X"af",X"4e",X"af",X"eb",X"4e",X"eb",X"4e",X"1c",X"10",X"3b",X"3b",X"74",X"3b",X"c7",X"c7",X"c7",X"c7",X"4c",X"00",X"00",X"f4",X"3c",X"8f",X"4f",X"fb",X"a4",X"a4",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"a4",X"8f",X"3c",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"9e",X"aa",X"7c",X"9e",X"98",X"0b",X"0b",X"1b",X"03",X"1a",X"1a",X"03",X"b2",X"03",X"19",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"27",X"19",X"71",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"75",X"b2",X"27",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"75",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"aa",X"2c",X"aa",X"33",X"1b",X"0b",X"1b",X"61",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"19",X"71",X"19",X"71",X"75",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"75",X"03",X"03",X"b2",X"27",X"1a",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"71",X"d8",X"2e",X"2e",X"1b",X"0b",X"0b",X"3c",X"39",X"d1",X"d1",X"d1",X"d1",X"57",X"d1",X"57",X"d1",X"39",X"39",X"4a",X"ae",X"39",X"ae",X"70",X"ae",X"82",X"82",X"ae",X"f3",X"22",X"f3",X"f3",X"f3",X"4e",X"3b",X"3b",X"8b",X"af",X"8b",X"af",X"2e",X"3b",X"1c",X"bb",X"bb",X"b9",X"b9",X"b9",X"b9",X"bb",X"c1",X"07",X"c1",X"bb",X"1c",X"10",X"10",X"1c",X"10",X"1c",X"3b",X"3b",X"4c",X"c7",X"3b",X"4c",X"c7",X"2e",X"c7",X"c7",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"f4",X"8f",X"a4",X"8f",X"a4",X"a4",X"8f",X"a4",X"a4",X"8f",X"a4",X"a4",X"8f",X"a4",X"3c",X"f4",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"aa",X"9e",X"aa",X"98",X"0b",X"1b",X"0b",X"19",X"03",X"03",X"03",X"19",X"03",X"b2",X"03",X"03",X"19",X"03",X"19",X"03",X"b2",X"27",X"75",X"71",X"03",X"19",X"03",X"b2",X"27",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"d8",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"71",X"19",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"3c",X"0b",X"0b",X"3b",X"6d",X"f0",X"3f",X"6d",
    X"aa",X"12",X"aa",X"aa",X"98",X"0b",X"0b",X"0b",X"2f",X"03",X"75",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"03",X"b2",X"27",X"19",X"03",X"19",X"03",X"71",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"03",X"14",X"09",X"2e",X"2e",X"1b",X"0b",X"0b",X"3c",X"39",X"d1",X"ff",X"d1",X"d1",X"d1",X"39",X"1f",X"d1",X"39",X"fb",X"82",X"39",X"ae",X"ae",X"ae",X"ae",X"f3",X"f3",X"f3",X"f3",X"22",X"af",X"8b",X"3b",X"8b",X"af",X"22",X"46",X"d7",X"2e",X"2e",X"3b",X"3b",X"1c",X"bb",X"07",X"9b",X"bb",X"07",X"c1",X"bb",X"bb",X"ce",X"10",X"1c",X"10",X"1c",X"10",X"3b",X"3b",X"4c",X"c7",X"74",X"3b",X"3b",X"4c",X"9a",X"2e",X"2e",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"fb",X"a4",X"8f",X"a4",X"a4",X"8f",X"a4",X"a4",X"8f",X"a4",X"8f",X"a4",X"8f",X"a4",X"3c",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"79",X"6d",X"f0",X"6d",X"aa",X"7c",X"aa",X"aa",X"33",X"0b",X"0b",X"0b",X"03",X"b2",X"27",X"19",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"19",X"b2",X"27",X"19",X"71",X"19",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"27",X"19",X"b2",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"19",X"0b",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"aa",X"7c",X"9e",X"98",X"0b",X"1b",X"0b",X"f0",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"27",X"1a",X"03",X"b2",X"03",X"b2",X"27",X"1a",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"03",X"71",X"d8",X"03",X"14",X"09",X"ec",X"2e",X"2e",X"2e",X"1b",X"0b",X"0b",X"3c",X"82",X"39",X"d1",X"ff",X"d1",X"39",X"d1",X"39",X"39",X"4a",X"ae",X"82",X"70",X"ae",X"f3",X"ae",X"f3",X"f3",X"22",X"8b",X"f3",X"4e",X"3b",X"4e",X"22",X"46",X"22",X"f3",X"46",X"4e",X"af",X"3b",X"3b",X"10",X"1c",X"bb",X"07",X"c1",X"bb",X"ce",X"10",X"1c",X"10",X"10",X"ce",X"3b",X"3b",X"3b",X"4c",X"c7",X"2e",X"74",X"4c",X"17",X"3b",X"4c",X"9a",X"2e",X"00",X"00",X"fb",X"00",X"a4",X"91",X"f4",X"fb",X"a4",X"8f",X"a4",X"8f",X"a4",X"8f",X"a4",X"8f",X"a4",X"8f",X"a4",X"3c",X"fb",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"9e",X"aa",X"9e",X"7c",X"61",X"0b",X"0b",X"1b",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"75",X"03",X"b2",X"03",X"03",X"19",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"b2",X"27",X"03",X"1a",X"03",X"1a",X"03",X"19",X"71",X"27",X"1a",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"19",X"b2",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"75",X"03",X"71",X"19",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"b2",X"03",X"19",X"71",X"1b",X"0b",X"0b",X"3b",X"f0",X"6d",X"3f",X"6d",
    X"aa",X"2c",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"79",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"1a",X"03",X"19",X"71",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"03",X"14",X"09",X"68",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"1b",X"0b",X"0b",X"3c",X"82",X"39",X"d1",X"ff",X"39",X"fb",X"39",X"ae",X"39",X"ae",X"82",X"ae",X"82",X"82",X"ae",X"f3",X"f3",X"f3",X"6f",X"8b",X"c6",X"af",X"2e",X"2e",X"d7",X"22",X"46",X"eb",X"8b",X"cd",X"3b",X"3b",X"3b",X"10",X"1c",X"10",X"10",X"1c",X"10",X"10",X"1c",X"3b",X"33",X"3b",X"4c",X"4c",X"c7",X"2e",X"74",X"4c",X"9a",X"03",X"3b",X"3b",X"3b",X"4c",X"00",X"00",X"f4",X"3c",X"8f",X"fb",X"f4",X"91",X"00",X"3c",X"3c",X"00",X"fb",X"fb",X"3c",X"3c",X"3c",X"3c",X"3c",X"fb",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"75",X"03",X"71",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"19",X"0b",X"1b",X"0b",X"98",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"12",X"aa",X"9e",X"98",X"1b",X"0b",X"0b",X"2f",X"03",X"b2",X"03",X"19",X"71",X"75",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"03",X"03",X"14",X"14",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"1b",X"0b",X"3c",X"0b",X"82",X"39",X"d1",X"39",X"d1",X"39",X"ae",X"82",X"39",X"ae",X"f3",X"ae",X"f3",X"82",X"f3",X"4e",X"f3",X"4e",X"3b",X"8b",X"2e",X"2e",X"d7",X"46",X"22",X"8b",X"af",X"3b",X"0b",X"2e",X"7f",X"58",X"3b",X"ad",X"1b",X"ad",X"3b",X"3b",X"3b",X"3b",X"2e",X"c7",X"4c",X"c7",X"2e",X"2e",X"74",X"4c",X"c7",X"03",X"b2",X"03",X"1b",X"3b",X"00",X"00",X"fb",X"00",X"a4",X"fb",X"fb",X"3c",X"a4",X"8f",X"a4",X"3c",X"f4",X"3c",X"8f",X"a4",X"a4",X"a4",X"a4",X"3c",X"91",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"3b",X"6d",X"f0",X"6d",X"f0",X"9e",X"aa",X"aa",X"92",X"61",X"0b",X"0b",X"0b",X"03",X"b2",X"27",X"03",X"1a",X"03",X"b2",X"27",X"75",X"71",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"b2",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"03",X"0b",X"0b",X"1b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"6d",X"aa",X"7c",X"61",X"0b",X"83",X"1b",X"ed",X"03",X"75",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"19",X"03",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"03",X"b2",X"03",X"71",X"d8",X"03",X"d8",X"14",X"ec",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"3c",X"0b",X"3c",X"0b",X"3c",X"82",X"39",X"ae",X"39",X"ae",X"82",X"70",X"ae",X"f3",X"ae",X"f3",X"22",X"f3",X"8b",X"f3",X"3b",X"3b",X"4e",X"22",X"46",X"22",X"8b",X"4e",X"17",X"cd",X"1b",X"0b",X"2e",X"1a",X"03",X"03",X"03",X"03",X"2e",X"2e",X"2e",X"2e",X"c7",X"c7",X"c7",X"2e",X"2e",X"74",X"4c",X"c7",X"2e",X"03",X"03",X"03",X"1a",X"03",X"00",X"00",X"f4",X"3c",X"a4",X"91",X"f4",X"a4",X"8f",X"a4",X"8f",X"3c",X"91",X"a4",X"a4",X"8f",X"a4",X"8f",X"8f",X"a4",X"3c",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"7c",X"aa",X"60",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"b2",X"03",X"03",X"19",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"03",X"75",X"03",X"b2",X"03",X"1a",X"03",X"75",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"d8",X"75",X"03",X"71",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"b2",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"9e",X"36",X"9e",X"aa",X"98",X"0b",X"1b",X"0b",X"79",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"06",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"75",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"b2",X"03",X"1a",X"03",X"b2",X"19",X"03",X"03",X"03",X"14",X"14",X"68",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"2e",X"2e",X"1b",X"0b",X"0b",X"00",X"0b",X"b8",X"ae",X"82",X"ae",X"ae",X"f3",X"ae",X"f3",X"f3",X"f3",X"48",X"f3",X"4e",X"8b",X"3b",X"3b",X"af",X"8b",X"af",X"af",X"3b",X"3b",X"0b",X"0b",X"3c",X"2e",X"03",X"03",X"b2",X"2e",X"2e",X"2e",X"2e",X"c7",X"c7",X"c7",X"2e",X"2e",X"2e",X"2e",X"74",X"4c",X"c7",X"2e",X"03",X"03",X"b2",X"19",X"b2",X"00",X"00",X"fb",X"00",X"8f",X"4f",X"fb",X"8f",X"a4",X"8f",X"a4",X"3c",X"4f",X"a4",X"8f",X"a4",X"8f",X"a4",X"a4",X"a4",X"3c",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"1b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"03",X"75",X"03",X"b2",X"03",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"d8",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"03",X"03",X"0b",X"0b",X"0b",X"3b",X"f0",X"6d",X"3f",X"6d",
    X"aa",X"60",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"2f",X"03",X"19",X"03",X"b2",X"27",X"1a",X"03",X"03",X"19",X"b2",X"27",X"19",X"03",X"75",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"03",X"b2",X"27",X"19",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"71",X"03",X"19",X"03",X"1a",X"03",X"03",X"03",X"03",X"d8",X"14",X"09",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"14",X"03",X"2e",X"2e",X"3c",X"0b",X"1b",X"0b",X"00",X"0b",X"82",X"ae",X"82",X"f3",X"ae",X"f3",X"22",X"f3",X"4e",X"f3",X"8b",X"af",X"3b",X"3b",X"3b",X"3b",X"3b",X"3b",X"3c",X"0b",X"3c",X"0b",X"30",X"03",X"1a",X"2e",X"2e",X"c7",X"c7",X"c7",X"c7",X"2e",X"2e",X"2e",X"2e",X"2e",X"4c",X"4c",X"c7",X"2e",X"d8",X"d8",X"03",X"03",X"03",X"03",X"00",X"00",X"f4",X"3c",X"a4",X"fb",X"f4",X"a4",X"3c",X"3c",X"3c",X"3c",X"3c",X"8f",X"3c",X"f4",X"3c",X"3c",X"3c",X"8f",X"3c",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"c6",X"6d",X"f0",X"6d",X"f0",X"aa",X"aa",X"7c",X"9e",X"61",X"0b",X"0b",X"1b",X"03",X"b2",X"03",X"03",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"75",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"75",X"03",X"03",X"b2",X"19",X"71",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"75",X"03",X"19",X"b2",X"19",X"3c",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"aa",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"61",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"71",X"19",X"71",X"19",X"71",X"03",X"03",X"14",X"ec",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"14",X"03",X"03",X"03",X"2e",X"2e",X"3c",X"0b",X"0b",X"0b",X"00",X"0b",X"eb",X"ae",X"f3",X"f3",X"f3",X"6f",X"f3",X"eb",X"4e",X"8b",X"4e",X"8b",X"4e",X"38",X"1b",X"0b",X"0b",X"3c",X"0b",X"0b",X"2e",X"03",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"4c",X"4c",X"c7",X"c7",X"2e",X"2e",X"03",X"03",X"03",X"03",X"b2",X"19",X"00",X"00",X"fb",X"00",X"8f",X"4f",X"fb",X"8f",X"a4",X"a4",X"8f",X"a4",X"8f",X"a4",X"3c",X"fb",X"8f",X"a4",X"8f",X"a4",X"3c",X"f4",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"6d",X"12",X"aa",X"aa",X"98",X"1b",X"83",X"0b",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"19",X"71",X"75",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"b2",X"03",X"75",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"03",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"f0",
    X"9e",X"7c",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"2f",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"27",X"19",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"03",X"03",X"03",X"14",X"09",X"68",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"09",X"a7",X"03",X"03",X"03",X"b2",X"03",X"2e",X"2e",X"1b",X"1b",X"0b",X"00",X"0b",X"1b",X"0b",X"00",X"eb",X"f3",X"8b",X"4e",X"8b",X"eb",X"8b",X"af",X"8b",X"4e",X"0b",X"0b",X"3c",X"0b",X"0b",X"3c",X"2e",X"03",X"1a",X"03",X"03",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"c7",X"c7",X"2e",X"2e",X"2e",X"14",X"03",X"03",X"b2",X"27",X"75",X"03",X"00",X"00",X"f4",X"3c",X"a4",X"fb",X"f4",X"a4",X"8f",X"a4",X"8f",X"a4",X"a4",X"8f",X"3c",X"fb",X"a4",X"8f",X"a4",X"8f",X"3c",X"fb",X"00",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"7c",X"9e",X"98",X"0b",X"1b",X"0b",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"03",X"75",X"03",X"b2",X"03",X"03",X"19",X"03",X"71",X"19",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"19",X"71",X"19",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"27",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"b2",X"19",X"03",X"b2",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"0b",X"0b",X"1b",X"17",X"6d",X"f0",X"6d",X"6d",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"1b",X"83",X"2f",X"03",X"19",X"71",X"19",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"b2",X"27",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"03",X"03",X"14",X"09",X"ec",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"14",X"14",X"03",X"71",X"03",X"19",X"03",X"b2",X"03",X"21",X"2e",X"2e",X"1b",X"0b",X"00",X"0b",X"0b",X"0b",X"00",X"0b",X"3c",X"eb",X"8b",X"4e",X"8b",X"4e",X"8b",X"3c",X"0b",X"00",X"0b",X"3c",X"0b",X"2e",X"27",X"19",X"71",X"03",X"14",X"09",X"a7",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"14",X"03",X"03",X"03",X"03",X"b2",X"03",X"03",X"00",X"00",X"fb",X"00",X"8f",X"fb",X"fb",X"f4",X"8f",X"a4",X"8f",X"a4",X"8f",X"3c",X"91",X"f4",X"8f",X"a4",X"a4",X"3c",X"f4",X"fb",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"f0",X"aa",X"60",X"aa",X"aa",X"98",X"0b",X"1b",X"0b",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"03",X"03",X"75",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"71",X"19",X"03",X"1a",X"03",X"19",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"1b",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"f0",
    X"aa",X"7c",X"aa",X"12",X"98",X"0b",X"0b",X"1b",X"ed",X"03",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"27",X"1a",X"03",X"19",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"19",X"71",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"03",X"03",X"03",X"14",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"14",X"03",X"03",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"1a",X"ec",X"2e",X"2e",X"1b",X"3c",X"1b",X"0b",X"3c",X"0b",X"0b",X"00",X"0b",X"3c",X"eb",X"af",X"0b",X"0b",X"0b",X"00",X"0b",X"2e",X"03",X"b2",X"27",X"03",X"03",X"03",X"14",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"14",X"d8",X"03",X"03",X"71",X"19",X"03",X"1a",X"00",X"00",X"f4",X"00",X"a4",X"91",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"91",X"f4",X"fb",X"f4",X"3c",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"9e",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"03",X"1a",X"03",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"19",X"b2",X"27",X"19",X"b2",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"27",X"75",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"0b",X"0b",X"0b",X"3b",X"3f",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"9e",X"aa",X"98",X"0b",X"1b",X"0b",X"79",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"71",X"d8",X"14",X"09",X"68",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"14",X"03",X"03",X"71",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"2e",X"2e",X"2e",X"2e",X"1b",X"0b",X"3c",X"0b",X"0b",X"0b",X"0b",X"0b",X"3c",X"0b",X"1b",X"0b",X"2e",X"03",X"1a",X"03",X"b2",X"03",X"03",X"d8",X"14",X"09",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"68",X"14",X"03",X"03",X"03",X"03",X"b2",X"03",X"00",X"00",X"fb",X"00",X"00",X"a4",X"4f",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"f4",X"fb",X"00",X"00",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"0b",X"3c",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"19",X"b2",X"27",X"19",X"71",X"03",X"03",X"b2",X"03",X"03",X"b2",X"27",X"19",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"d8",X"19",X"71",X"19",X"03",X"19",X"03",X"1a",X"03",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"19",X"03",X"75",X"03",X"b2",X"03",X"19",X"03",X"03",X"19",X"b2",X"27",X"19",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"b2",X"03",X"75",X"03",X"0b",X"00",X"0b",X"98",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"60",X"98",X"1b",X"0b",X"0b",X"2f",X"03",X"b2",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"75",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"03",X"75",X"03",X"b2",X"03",X"03",X"19",X"03",X"14",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"14",X"03",X"27",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"19",X"ec",X"2e",X"2e",X"1b",X"0b",X"3c",X"0b",X"3c",X"0b",X"0b",X"ec",X"2e",X"03",X"b2",X"03",X"19",X"03",X"03",X"03",X"14",X"14",X"ec",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"09",X"14",X"03",X"03",X"03",X"1a",X"03",X"03",X"00",X"00",X"f4",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"f4",X"fb",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"cd",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"9e",X"aa",X"9e",X"98",X"0b",X"1b",X"0b",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"b2",X"27",X"75",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"19",X"71",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"b2",X"19",X"03",X"b2",X"03",X"19",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"75",X"03",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"0b",X"0b",X"0b",X"3b",X"f0",X"6d",X"f0",X"6d",
    X"aa",X"9e",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"61",X"03",X"75",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"19",X"71",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"19",X"71",X"19",X"71",X"19",X"71",X"19",X"03",X"1a",X"03",X"71",X"d8",X"d8",X"14",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"09",X"14",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"b2",X"27",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"71",X"30",X"2e",X"2e",X"ec",X"0b",X"1b",X"2e",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"71",X"14",X"14",X"68",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"14",X"03",X"03",X"b2",X"27",X"19",X"1a",X"00",X"00",X"00",X"f4",X"fb",X"f4",X"f4",X"fb",X"f4",X"f4",X"fb",X"f4",X"f4",X"fb",X"f4",X"fb",X"f4",X"f4",X"fb",X"f4",X"f4",X"fb",X"f4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",X"7c",X"0d",X"7c",X"aa",X"ba",X"0b",X"0b",X"0b",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"75",X"03",X"1a",X"03",X"75",X"03",X"b2",X"03",X"1a",X"03",X"1a",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"71",X"19",X"03",X"b2",X"19",X"03",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"19",X"03",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"1a",X"03",X"19",X"03",X"03",X"b2",X"19",X"03",X"b2",X"03",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"71",X"19",X"03",X"1a",X"03",X"71",X"19",X"71",X"27",X"1a",X"03",X"19",X"03",X"19",X"03",X"03",X"1a",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"0b",X"0b",X"1b",X"33",X"6d",X"f0",X"6d",X"3f",
    X"aa",X"7c",X"0d",X"9e",X"98",X"0b",X"1b",X"0b",X"2f",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"1a",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"b2",X"03",X"75",X"03",X"03",X"75",X"03",X"03",X"b2",X"03",X"03",X"03",X"03",X"14",X"09",X"68",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"14",X"03",X"03",X"03",X"03",X"1a",X"03",X"b2",X"27",X"03",X"b2",X"03",X"19",X"b2",X"27",X"19",X"1a",X"03",X"b2",X"27",X"19",X"03",X"03",X"b2",X"19",X"2e",X"30",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"03",X"03",X"14",X"14",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"14",X"03",X"03",X"03",X"b2",X"03",X"03",X"00",X"00",X"00",X"3c",X"00",X"00",X"00",X"3c",X"00",X"3c",X"00",X"3c",X"00",X"3c",X"00",X"00",X"00",X"3c",X"00",X"3c",X"00",X"3c",X"00",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"6d",X"f0",X"6d",X"3f",X"aa",X"2c",X"aa",X"9e",X"54",X"0b",X"0b",X"1b",X"03",X"b2",X"19",X"71",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"03",X"19",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"19",X"71",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"19",X"71",X"27",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"19",X"71",X"19",X"03",X"71",X"19",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"19",X"71",X"27",X"1a",X"03",X"b2",X"03",X"1a",X"1b",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"7c",X"aa",X"61",X"0b",X"0b",X"0b",X"79",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"1a",X"03",X"03",X"b2",X"19",X"03",X"03",X"b2",X"03",X"19",X"03",X"1a",X"03",X"b2",X"03",X"75",X"03",X"03",X"b2",X"19",X"71",X"03",X"1a",X"03",X"19",X"03",X"71",X"03",X"d8",X"14",X"09",X"ec",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"14",X"27",X"03",X"b2",X"19",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"b2",X"03",X"03",X"1a",X"03",X"b2",X"03",X"03",X"d8",X"14",X"09",X"ec",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"14",X"27",X"03",X"71",X"19",X"03",X"b2",X"00",X"00",X"00",X"70",X"3c",X"f3",X"3c",X"82",X"3c",X"82",X"3c",X"70",X"3c",X"82",X"3c",X"f3",X"3c",X"82",X"3c",X"82",X"3c",X"70",X"3c",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"12",X"aa",X"aa",X"84",X"0b",X"1b",X"0b",X"19",X"03",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"03",X"19",X"b2",X"19",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"1a",X"03",X"03",X"19",X"b2",X"27",X"19",X"03",X"19",X"b2",X"19",X"03",X"19",X"03",X"19",X"03",X"75",X"03",X"03",X"19",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"1a",X"03",X"1a",X"03",X"03",X"1a",X"03",X"b2",X"27",X"19",X"03",X"19",X"03",X"75",X"03",X"03",X"19",X"03",X"1a",X"03",X"19",X"71",X"19",X"03",X"1a",X"03",X"b2",X"03",X"19",X"03",X"19",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"03",X"1b",X"0b",X"0b",X"53",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"9e",X"aa",X"60",X"98",X"0b",X"1b",X"83",X"2f",X"27",X"b2",X"03",X"19",X"03",X"b2",X"27",X"19",X"03",X"b2",X"27",X"19",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"b2",X"27",X"19",X"03",X"b2",X"27",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"b2",X"03",X"03",X"03",X"14",X"14",X"14",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"09",X"14",X"d8",X"03",X"03",X"03",X"03",X"1a",X"03",X"19",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"1a",X"03",X"03",X"19",X"03",X"03",X"14",X"09",X"09",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"2e",X"ec",X"09",X"14",X"d8",X"03",X"03",X"03",X"1a",X"03",X"00",X"00",X"00",X"82",X"3c",X"70",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"70",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"3c",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"6d",X"aa",X"9e",X"aa",X"7c",X"61",X"0b",X"0b",X"1b",X"03",X"b2",X"19",X"71",X"19",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"b2",X"03",X"1a",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"19",X"71",X"19",X"71",X"19",X"71",X"19",X"03",X"71",X"19",X"71",X"19",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"19",X"71",X"19",X"71",X"19",X"71",X"19",X"03",X"71",X"19",X"71",X"19",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"19",X"71",X"19",X"71",X"19",X"71",X"19",X"03",X"71",X"19",X"71",X"19",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"03",X"b2",X"19",X"71",X"19",X"71",X"19",X"b2",X"83",X"0b",X"0b",X"33",X"6d",X"3f",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"aa",X"ba",X"0b",X"0b",X"1b",X"53",X"79",X"79",X"79",X"2f",X"79",X"79",X"2f",X"79",X"79",X"79",X"ed",X"f0",X"77",X"79",X"79",X"2f",X"79",X"2f",X"79",X"2f",X"79",X"79",X"2f",X"79",X"79",X"79",X"79",X"77",X"79",X"2f",X"79",X"79",X"ed",X"79",X"2f",X"79",X"2f",X"79",X"77",X"f0",X"77",X"2f",X"f0",X"77",X"79",X"79",X"79",X"77",X"f0",X"f0",X"79",X"3f",X"63",X"20",X"16",X"16",X"69",X"16",X"69",X"16",X"b1",X"16",X"16",X"20",X"3f",X"28",X"28",X"79",X"61",X"2f",X"79",X"79",X"2f",X"79",X"2f",X"79",X"2f",X"79",X"79",X"2f",X"79",X"2f",X"79",X"2f",X"79",X"79",X"79",X"77",X"f0",X"77",X"79",X"2f",X"79",X"79",X"2f",X"79",X"2f",X"28",X"79",X"f0",X"0d",X"63",X"63",X"69",X"16",X"b1",X"16",X"b1",X"16",X"16",X"b1",X"63",X"3f",X"28",X"79",X"f0",X"77",X"2f",X"79",X"79",X"00",X"00",X"00",X"82",X"00",X"82",X"00",X"82",X"00",X"82",X"00",X"82",X"00",X"82",X"00",X"82",X"00",X"82",X"00",X"82",X"00",X"82",X"00",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0b",X"0b",X"33",X"6d",X"3f",X"6d",X"f0",X"7c",X"aa",X"6d",X"aa",X"84",X"0b",X"1b",X"0b",X"19",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"1a",X"03",X"19",X"03",X"75",X"03",X"19",X"03",X"19",X"03",X"19",X"03",X"75",X"03",X"19",X"03",X"75",X"03",X"75",X"03",X"19",X"03",X"75",X"03",X"75",X"03",X"19",X"03",X"19",X"03",X"19",X"03",X"75",X"03",X"19",X"03",X"75",X"03",X"75",X"03",X"19",X"03",X"75",X"03",X"75",X"03",X"19",X"03",X"19",X"03",X"19",X"03",X"75",X"03",X"19",X"03",X"75",X"03",X"75",X"03",X"19",X"03",X"75",X"03",X"75",X"03",X"19",X"03",X"19",X"03",X"19",X"03",X"75",X"03",X"19",X"03",X"75",X"03",X"75",X"03",X"19",X"03",X"75",X"03",X"75",X"03",X"19",X"03",X"19",X"03",X"19",X"03",X"75",X"03",X"19",X"03",X"0b",X"3c",X"0b",X"17",X"f0",X"6d",X"f0",X"6d",
    X"9e",X"aa",X"9e",X"2c",X"61",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"1b",X"0b",X"1b",X"0b",X"1b",X"1b",X"0b",X"1b",X"0b",X"83",X"0b",X"1b",X"83",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"0b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"0b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"0b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"0b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"0b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"0b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"0b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"83",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"83",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"83",X"0b",X"1b",X"0b",X"1b",X"83",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"1b",X"83",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"0b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"0b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"0b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"0b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"0b",X"1b",X"0b",X"3b",X"f0",X"6d",X"f0",X"6d",X"aa",X"aa",X"12",X"aa",X"98",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"83",X"0b",X"0b",X"1b",X"83",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"0b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"0b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"0b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"0b",X"83",X"0b",X"1b",X"0b",X"83",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"1b",X"0b",X"1b",X"1b",X"0b",X"83",X"1b",X"33",X"6d",X"f0",X"6d",X"f0",
    X"aa",X"7c",X"aa",X"aa",X"98",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"33",X"6d",X"f0",X"54",X"3f",X"aa",X"60",X"aa",X"7c",X"61",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"33",X"f0",X"6d",X"f0",X"3f",
    X"aa",X"9e",X"aa",X"92",X"61",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"ad",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"ad",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"33",X"f0",X"6d",X"3f",X"6d",X"aa",X"aa",X"9e",X"aa",X"98",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"0b",X"1b",X"0b",X"1b",X"0b",X"0b",X"0b",X"33",X"6d",X"3f",X"54",X"6d",
    X"aa",X"7c",X"aa",X"ba",X"3b",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"84",X"98",X"ba",X"98",X"98",X"33",X"61",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"33",X"98",X"98",X"ba",X"98",X"33",X"98",X"61",X"98",X"98",X"98",X"ba",X"98",X"84",X"98",X"98",X"61",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"33",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"84",X"98",X"98",X"98",X"33",X"98",X"98",X"98",X"ba",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"17",X"61",X"6d",X"f0",X"6d",X"9e",X"7c",X"aa",X"98",X"33",X"54",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"98",X"98",X"61",X"98",X"98",X"33",X"98",X"84",X"61",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"61",X"98",X"17",X"98",X"f0",X"6d",X"3f",
    X"9e",X"aa",X"98",X"17",X"6d",X"aa",X"9e",X"aa",X"aa",X"12",X"2c",X"aa",X"aa",X"12",X"2c",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"aa",X"2c",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"60",X"aa",X"92",X"aa",X"aa",X"7c",X"aa",X"7c",X"aa",X"aa",X"2c",X"42",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"2c",X"aa",X"42",X"6d",X"aa",X"7c",X"aa",X"92",X"aa",X"60",X"aa",X"7c",X"9e",X"aa",X"7c",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"aa",X"9e",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"60",X"aa",X"2c",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"61",X"17",X"98",X"6d",X"f0",X"aa",X"aa",X"98",X"33",X"98",X"12",X"2c",X"aa",X"9e",X"aa",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"0d",X"9e",X"7c",X"aa",X"aa",X"7c",X"9e",X"aa",X"aa",X"12",X"aa",X"9e",X"60",X"aa",X"aa",X"7c",X"aa",X"74",X"17",X"98",X"6d",X"f0",
    X"aa",X"74",X"17",X"ba",X"aa",X"7c",X"0d",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"aa",X"aa",X"aa",X"aa",X"60",X"aa",X"9e",X"aa",X"aa",X"aa",X"12",X"aa",X"6d",X"aa",X"9e",X"aa",X"aa",X"aa",X"12",X"aa",X"6d",X"aa",X"9e",X"aa",X"9e",X"aa",X"aa",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"9e",X"aa",X"aa",X"7c",X"0d",X"60",X"aa",X"7c",X"aa",X"aa",X"9e",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"9e",X"aa",X"9e",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"ba",X"17",X"33",X"f0",X"7c",X"ba",X"33",X"98",X"aa",X"aa",X"9e",X"aa",X"7c",X"0d",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"aa",X"60",X"aa",X"aa",X"aa",X"98",X"3b",X"98",X"54",
    X"98",X"3b",X"6d",X"aa",X"60",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"12",X"2c",X"aa",X"92",X"aa",X"7c",X"aa",X"aa",X"12",X"2c",X"aa",X"92",X"aa",X"7c",X"aa",X"aa",X"12",X"2c",X"aa",X"92",X"aa",X"7c",X"aa",X"aa",X"7c",X"aa",X"60",X"aa",X"7c",X"aa",X"6d",X"36",X"6d",X"aa",X"7c",X"aa",X"60",X"aa",X"7c",X"aa",X"aa",X"12",X"aa",X"7c",X"aa",X"7c",X"aa",X"9e",X"aa",X"9e",X"aa",X"7c",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"98",X"3b",X"0b",X"ba",X"17",X"98",X"aa",X"92",X"aa",X"7c",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"aa",X"9e",X"aa",X"7c",X"9e",X"aa",X"7c",X"9e",X"7c",X"aa",X"6d",X"3b",X"33",
    X"0b",X"61",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"0d",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"60",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"60",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"60",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"60",X"aa",X"9e",X"aa",X"9e",X"aa",X"9e",X"aa",X"9e",X"aa",X"9e",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"60",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"98",X"0b",X"61",X"98",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"7c",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"aa",X"9e",X"aa",X"98",X"0b", others=>"00");
end package;