library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.graphics_pkg.all;

package sprite_pkg is
    constant TRANSPARENT_PIXEL : pixel_type := X"01";
end;