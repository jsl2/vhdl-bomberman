use work.graphics_pkg.all;

package powerup_pkg is    
    type powerup_rom_type is array(0 to (2**11 - 1)) of pixel_type;    
    
    constant POWERUP_SPRITES : powerup_rom_type := 
   (X"48",X"48",X"6f",X"48",X"48",X"6f",X"48",X"48",X"6f",X"48",X"6f",X"48",X"48",X"6f",X"48",X"6f",
    X"6f",X"4b",X"4b",X"4b",X"4b",X"00",X"00",X"00",X"3c",X"00",X"3c",X"4b",X"00",X"3c",X"4b",X"48",
    X"48",X"4b",X"4b",X"00",X"00",X"23",X"23",X"23",X"00",X"23",X"12",X"00",X"4b",X"46",X"00",X"48",
    X"6f",X"4b",X"00",X"23",X"23",X"23",X"23",X"00",X"12",X"2e",X"00",X"4b",X"00",X"00",X"4b",X"6f",
    X"48",X"4b",X"00",X"23",X"12",X"12",X"12",X"00",X"12",X"4b",X"00",X"00",X"23",X"00",X"4b",X"48",
    X"6f",X"00",X"23",X"12",X"12",X"2e",X"12",X"00",X"23",X"12",X"4b",X"12",X"23",X"00",X"00",X"48",
    X"48",X"00",X"23",X"12",X"12",X"12",X"12",X"12",X"00",X"23",X"12",X"23",X"00",X"00",X"00",X"6f",
    X"6f",X"3c",X"ba",X"12",X"12",X"12",X"12",X"12",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"48",
    X"48",X"00",X"23",X"12",X"12",X"12",X"12",X"12",X"23",X"23",X"23",X"00",X"00",X"00",X"00",X"48",
    X"6f",X"00",X"23",X"23",X"12",X"12",X"12",X"23",X"23",X"23",X"00",X"00",X"00",X"00",X"00",X"6f",
    X"48",X"00",X"00",X"23",X"23",X"23",X"23",X"23",X"23",X"ba",X"00",X"00",X"00",X"00",X"00",X"48",
    X"6f",X"4b",X"00",X"23",X"23",X"23",X"23",X"23",X"23",X"3c",X"00",X"00",X"00",X"00",X"4b",X"48",
    X"48",X"4b",X"00",X"00",X"23",X"23",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4b",X"6f",
    X"6f",X"4b",X"4b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4b",X"4b",X"48",
    X"48",X"4b",X"4b",X"4b",X"4b",X"00",X"00",X"3c",X"00",X"00",X"00",X"4b",X"4b",X"4b",X"4b",X"6f",
    X"6f",X"48",X"48",X"6f",X"48",X"48",X"6f",X"48",X"48",X"6f",X"48",X"48",X"6f",X"48",X"48",X"48",
    X"48",X"48",X"6f",X"48",X"48",X"6f",X"48",X"6f",X"48",X"48",X"6f",X"48",X"6f",X"48",X"48",X"6f",
    X"6f",X"4b",X"4b",X"4b",X"4b",X"4b",X"4b",X"cb",X"4b",X"4b",X"cb",X"4b",X"4b",X"cb",X"4b",X"f3",
    X"48",X"4b",X"4b",X"4b",X"4b",X"4b",X"cb",X"46",X"cb",X"cb",X"4f",X"cb",X"cb",X"46",X"cb",X"8b",
    X"6f",X"4b",X"4b",X"4b",X"cb",X"cb",X"46",X"4f",X"cb",X"4f",X"4f",X"cb",X"4f",X"46",X"cb",X"f3",
    X"48",X"4b",X"4b",X"cb",X"46",X"2e",X"2e",X"4f",X"4f",X"4f",X"4f",X"4f",X"4f",X"46",X"cb",X"48",
    X"6f",X"4b",X"cb",X"46",X"2e",X"2e",X"4f",X"4f",X"2e",X"4f",X"4f",X"4f",X"4f",X"46",X"cb",X"6f",
    X"48",X"4b",X"cb",X"2e",X"4f",X"00",X"2e",X"4f",X"00",X"2e",X"4f",X"4f",X"4f",X"46",X"cb",X"f3",
    X"6f",X"cb",X"46",X"4f",X"4f",X"00",X"2e",X"4f",X"00",X"2e",X"4f",X"4f",X"4f",X"46",X"cb",X"8b",
    X"48",X"cb",X"4f",X"4f",X"4f",X"00",X"2e",X"4f",X"00",X"2e",X"4f",X"4f",X"4f",X"46",X"cb",X"f3",
    X"6f",X"cb",X"4f",X"4f",X"2e",X"4f",X"4f",X"4f",X"4f",X"4f",X"4f",X"4f",X"4f",X"46",X"cb",X"48",
    X"48",X"cb",X"46",X"4f",X"cb",X"3c",X"00",X"00",X"00",X"00",X"4f",X"4f",X"46",X"cb",X"4b",X"6f",
    X"6f",X"cb",X"46",X"4f",X"4f",X"cb",X"8b",X"8b",X"00",X"46",X"4f",X"4f",X"46",X"67",X"4b",X"48",
    X"48",X"4b",X"cb",X"46",X"4f",X"4f",X"cb",X"cb",X"46",X"4f",X"4f",X"46",X"cb",X"4b",X"4b",X"8b",
    X"6f",X"4b",X"4b",X"cb",X"cb",X"4f",X"4f",X"4f",X"4f",X"46",X"cb",X"cb",X"7b",X"4b",X"4b",X"f3",
    X"48",X"4b",X"4b",X"4b",X"7b",X"cb",X"cb",X"cb",X"cb",X"cb",X"4b",X"4b",X"4b",X"4b",X"4b",X"8b",
    X"6f",X"48",X"48",X"6f",X"48",X"6f",X"48",X"48",X"6f",X"48",X"48",X"48",X"6f",X"48",X"48",X"6f",
    X"48",X"48",X"6f",X"48",X"48",X"6f",X"48",X"48",X"6f",X"48",X"6f",X"48",X"48",X"6f",X"48",X"48",
    X"6f",X"4b",X"4b",X"4b",X"4b",X"4b",X"00",X"cb",X"cb",X"cb",X"cb",X"cb",X"cb",X"00",X"4b",X"6f",
    X"48",X"4b",X"4b",X"4b",X"4b",X"4b",X"00",X"12",X"12",X"4b",X"2e",X"4b",X"12",X"00",X"4b",X"f3",
    X"6f",X"4b",X"4b",X"4b",X"4b",X"00",X"4f",X"4f",X"46",X"8b",X"2e",X"4b",X"12",X"00",X"4b",X"48",
    X"48",X"4b",X"4b",X"4b",X"4b",X"4b",X"00",X"12",X"12",X"4b",X"2e",X"4b",X"12",X"00",X"4b",X"6f",
    X"6f",X"4b",X"4b",X"4b",X"4b",X"00",X"4f",X"4f",X"46",X"8b",X"2e",X"4b",X"12",X"00",X"4b",X"48",
    X"48",X"4b",X"4b",X"00",X"00",X"00",X"00",X"12",X"12",X"4b",X"2e",X"4b",X"12",X"00",X"4b",X"f3",
    X"6f",X"4b",X"00",X"12",X"4b",X"4b",X"4b",X"4b",X"4b",X"4b",X"4b",X"4b",X"12",X"00",X"4b",X"48",
    X"48",X"00",X"12",X"4b",X"12",X"12",X"4b",X"4b",X"4b",X"4b",X"12",X"12",X"4b",X"12",X"00",X"6f",
    X"6f",X"3c",X"12",X"12",X"00",X"00",X"12",X"12",X"4b",X"12",X"00",X"00",X"12",X"12",X"00",X"f3",
    X"48",X"00",X"12",X"00",X"4f",X"4f",X"00",X"12",X"12",X"00",X"4f",X"4f",X"00",X"12",X"00",X"8b",
    X"6f",X"4b",X"00",X"4f",X"23",X"23",X"4f",X"00",X"00",X"4f",X"23",X"23",X"4f",X"00",X"00",X"f3",
    X"48",X"4b",X"00",X"46",X"23",X"23",X"fb",X"00",X"00",X"46",X"23",X"23",X"4f",X"00",X"4b",X"48",
    X"6f",X"4b",X"4b",X"00",X"46",X"fb",X"00",X"4b",X"4b",X"00",X"46",X"fb",X"00",X"4b",X"4b",X"6f",
    X"48",X"4b",X"4b",X"4b",X"3c",X"00",X"4b",X"4b",X"4b",X"4b",X"3c",X"00",X"4b",X"4b",X"4b",X"48",
    X"6f",X"48",X"48",X"6f",X"48",X"48",X"6f",X"48",X"48",X"6f",X"48",X"6f",X"48",X"48",X"6f",X"f3",
    X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",
    X"27",X"a0",X"a0",X"4b",X"a0",X"3c",X"3c",X"3c",X"3c",X"3c",X"3c",X"a0",X"3c",X"3c",X"a0",X"27",
    X"27",X"a0",X"4b",X"3c",X"00",X"74",X"ba",X"74",X"00",X"23",X"12",X"00",X"4b",X"46",X"3c",X"27",
    X"27",X"a0",X"3c",X"23",X"23",X"23",X"23",X"00",X"12",X"2e",X"00",X"4b",X"00",X"00",X"4b",X"27",
    X"27",X"a0",X"00",X"23",X"12",X"12",X"12",X"00",X"12",X"4b",X"00",X"00",X"23",X"00",X"4b",X"27",
    X"27",X"3c",X"74",X"12",X"12",X"2e",X"12",X"00",X"23",X"12",X"4b",X"12",X"23",X"00",X"00",X"27",
    X"27",X"3c",X"23",X"12",X"12",X"12",X"12",X"12",X"00",X"23",X"12",X"23",X"00",X"00",X"00",X"27",
    X"27",X"3c",X"74",X"12",X"12",X"12",X"12",X"12",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"27",
    X"27",X"3c",X"ba",X"12",X"12",X"12",X"12",X"12",X"23",X"23",X"23",X"00",X"00",X"00",X"00",X"27",
    X"27",X"3c",X"74",X"23",X"12",X"12",X"12",X"ba",X"23",X"ba",X"00",X"00",X"00",X"00",X"00",X"27",
    X"27",X"3c",X"00",X"23",X"23",X"ba",X"23",X"74",X"23",X"74",X"00",X"00",X"00",X"00",X"00",X"27",
    X"27",X"a0",X"3c",X"23",X"23",X"74",X"23",X"ba",X"23",X"3c",X"00",X"00",X"00",X"00",X"4b",X"27",
    X"27",X"a0",X"00",X"00",X"23",X"23",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4b",X"27",
    X"27",X"a0",X"4b",X"3c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4b",X"4b",X"27",
    X"27",X"a0",X"4b",X"4b",X"4b",X"00",X"00",X"3c",X"00",X"3c",X"00",X"a0",X"4b",X"a0",X"4b",X"27",
    X"27",X"27",X"36",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",
    X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",
    X"27",X"a0",X"a0",X"4b",X"a0",X"4b",X"a0",X"55",X"a0",X"a0",X"55",X"4b",X"a0",X"55",X"a0",X"27",
    X"27",X"a0",X"4b",X"4b",X"4b",X"4b",X"55",X"46",X"cb",X"cb",X"4f",X"cb",X"cb",X"46",X"cb",X"27",
    X"27",X"a0",X"4b",X"4b",X"55",X"cb",X"46",X"4f",X"cb",X"4f",X"4f",X"cb",X"4f",X"46",X"cb",X"27",
    X"27",X"a0",X"4b",X"cb",X"46",X"2e",X"2e",X"4f",X"4f",X"4f",X"4f",X"4f",X"4f",X"46",X"cb",X"27",
    X"27",X"a0",X"55",X"46",X"2e",X"2e",X"4f",X"4f",X"2e",X"4f",X"4f",X"4f",X"4f",X"46",X"cb",X"27",
    X"27",X"a0",X"cb",X"2e",X"4f",X"00",X"2e",X"4f",X"00",X"2e",X"4f",X"4f",X"4f",X"46",X"cb",X"27",
    X"27",X"bd",X"46",X"4f",X"4f",X"00",X"2e",X"4f",X"00",X"2e",X"4f",X"4f",X"4f",X"46",X"cb",X"27",
    X"27",X"55",X"fb",X"4f",X"4f",X"00",X"2e",X"4f",X"00",X"2e",X"4f",X"4f",X"4f",X"46",X"cb",X"27",
    X"27",X"55",X"4f",X"4f",X"2e",X"4f",X"4f",X"4f",X"4f",X"4f",X"4f",X"4f",X"4f",X"46",X"cb",X"27",
    X"27",X"55",X"46",X"4f",X"cb",X"00",X"00",X"00",X"00",X"00",X"fb",X"4f",X"46",X"cb",X"4b",X"27",
    X"27",X"55",X"46",X"4f",X"4f",X"cb",X"8b",X"8b",X"00",X"46",X"4f",X"4f",X"46",X"cb",X"4b",X"27",
    X"27",X"a0",X"cb",X"46",X"4f",X"4f",X"cb",X"cb",X"46",X"fb",X"4f",X"46",X"cb",X"4b",X"4b",X"27",
    X"27",X"a0",X"4b",X"cb",X"cb",X"4f",X"4f",X"4f",X"4f",X"46",X"cb",X"cb",X"4b",X"4b",X"4b",X"27",
    X"27",X"a0",X"4b",X"4b",X"4b",X"55",X"cb",X"cb",X"cb",X"cb",X"a0",X"4b",X"4b",X"4b",X"4b",X"27",
    X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",
    X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",
    X"27",X"a0",X"a0",X"4b",X"a0",X"4b",X"3c",X"bd",X"55",X"55",X"cb",X"55",X"55",X"3c",X"a0",X"27",
    X"27",X"a0",X"4b",X"4b",X"4b",X"4b",X"3c",X"12",X"12",X"4b",X"2e",X"4b",X"12",X"00",X"4b",X"27",
    X"27",X"a0",X"4b",X"4b",X"4b",X"3c",X"fb",X"4f",X"46",X"8b",X"2e",X"4b",X"12",X"00",X"4b",X"27",
    X"27",X"a0",X"4b",X"4b",X"4b",X"4b",X"00",X"12",X"12",X"4b",X"2e",X"4b",X"12",X"00",X"4b",X"27",
    X"27",X"a0",X"4b",X"4b",X"4b",X"3c",X"4f",X"4f",X"46",X"8b",X"2e",X"4b",X"12",X"00",X"a0",X"27",
    X"27",X"a0",X"4b",X"3c",X"00",X"00",X"00",X"12",X"12",X"4b",X"2e",X"4b",X"12",X"00",X"4b",X"27",
    X"27",X"a0",X"3c",X"12",X"4b",X"4b",X"4b",X"4b",X"4b",X"4b",X"4b",X"4b",X"12",X"00",X"4b",X"27",
    X"27",X"3c",X"12",X"4b",X"12",X"12",X"4b",X"4b",X"4b",X"4b",X"12",X"12",X"4b",X"12",X"00",X"27",
    X"27",X"3c",X"12",X"12",X"00",X"00",X"12",X"12",X"4b",X"12",X"00",X"00",X"12",X"12",X"00",X"27",
    X"27",X"3c",X"12",X"3c",X"4f",X"4f",X"00",X"12",X"12",X"00",X"4f",X"4f",X"00",X"12",X"00",X"27",
    X"27",X"a0",X"3c",X"fb",X"23",X"23",X"4f",X"00",X"00",X"4f",X"23",X"23",X"4f",X"00",X"00",X"27",
    X"27",X"a0",X"00",X"46",X"23",X"23",X"4f",X"00",X"00",X"46",X"23",X"23",X"4f",X"00",X"4b",X"27",
    X"27",X"a0",X"4b",X"00",X"46",X"4f",X"00",X"4b",X"4b",X"00",X"46",X"4f",X"00",X"4b",X"4b",X"27",
    X"27",X"a0",X"4b",X"4b",X"00",X"3c",X"4b",X"4b",X"4b",X"a0",X"00",X"3c",X"4b",X"4b",X"4b",X"27",
    X"27",X"27",X"36",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"36",others=>X"01"
    );
end package;