use work.graphics_pkg.all;

package bombs_pkg is
    constant MAX_BOMBS : integer := 9;
    constant MAX_BLAST_RADIUS : integer := 9;        
    
    constant small_bomb : bitmap_type := 
       ((X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"2e",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"2e",X"2e",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"00",X"00",X"53",X"ba",X"8c",X"8c",X"00",X"8c",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"00",X"53",X"ba",X"ba",X"53",X"2e",X"00",X"8c",X"00",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"00",X"9e",X"2e",X"9e",X"53",X"2e",X"00",X"00",X"8c",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"00",X"9e",X"9e",X"9e",X"9e",X"53",X"8c",X"8c",X"8c",X"8c",X"00",X"00",X"01",X"01"),
        (X"01",X"01",X"00",X"9e",X"2e",X"9e",X"9e",X"9e",X"53",X"8c",X"8c",X"53",X"53",X"00",X"01",X"01"),
        (X"01",X"01",X"00",X"9e",X"2e",X"9e",X"9e",X"9e",X"9e",X"53",X"53",X"53",X"53",X"00",X"01",X"01"),
        (X"01",X"01",X"00",X"9e",X"9e",X"9e",X"9e",X"9e",X"ba",X"ba",X"ba",X"53",X"53",X"00",X"01",X"01"),
        (X"01",X"01",X"00",X"ba",X"9e",X"9e",X"9e",X"ba",X"ba",X"ba",X"ba",X"53",X"53",X"00",X"01",X"01"),
        (X"01",X"01",X"01",X"00",X"ba",X"ba",X"ba",X"ba",X"ba",X"ba",X"53",X"53",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"00",X"53",X"53",X"ba",X"ba",X"ba",X"53",X"53",X"53",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"00",X"00",X"53",X"53",X"53",X"53",X"00",X"00",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"));
    
    constant medium_bomb : bitmap_type := 
       ((X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"2e",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"2e",X"2e",X"01"),
        (X"01",X"01",X"01",X"00",X"00",X"ba",X"ba",X"ba",X"ba",X"8c",X"8c",X"00",X"8c",X"00",X"01",X"01"),
        (X"01",X"01",X"00",X"ba",X"9e",X"2e",X"9e",X"ba",X"53",X"2e",X"00",X"8c",X"00",X"00",X"01",X"01"),
        (X"01",X"01",X"00",X"9e",X"9e",X"9e",X"9e",X"9e",X"53",X"2e",X"00",X"00",X"8c",X"00",X"01",X"01"),
        (X"01",X"00",X"9e",X"2e",X"2e",X"9e",X"9e",X"9e",X"53",X"8c",X"8c",X"8c",X"8c",X"53",X"00",X"01"),
        (X"01",X"00",X"9e",X"2e",X"2e",X"9e",X"9e",X"9e",X"9e",X"53",X"8c",X"8c",X"53",X"53",X"00",X"01"),
        (X"01",X"00",X"9e",X"9e",X"9e",X"9e",X"9e",X"9e",X"9e",X"ba",X"53",X"53",X"53",X"53",X"00",X"01"),
        (X"01",X"00",X"9e",X"9e",X"9e",X"9e",X"9e",X"9e",X"9e",X"ba",X"ba",X"53",X"53",X"53",X"00",X"01"),
        (X"01",X"00",X"9e",X"9e",X"9e",X"9e",X"9e",X"9e",X"ba",X"ba",X"ba",X"53",X"53",X"53",X"00",X"01"),
        (X"01",X"00",X"ba",X"9e",X"9e",X"9e",X"9e",X"ba",X"ba",X"ba",X"53",X"53",X"53",X"53",X"00",X"01"),
        (X"01",X"01",X"00",X"ba",X"ba",X"ba",X"ba",X"ba",X"ba",X"ba",X"53",X"53",X"53",X"00",X"01",X"01"),
        (X"01",X"01",X"00",X"53",X"ba",X"ba",X"ba",X"ba",X"53",X"53",X"53",X"53",X"53",X"00",X"01",X"01"),
        (X"01",X"01",X"01",X"00",X"00",X"53",X"53",X"53",X"53",X"53",X"53",X"00",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01"));
    
    constant large_bomb : bitmap_type := 
       ((X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"2e",X"2e",X"01"),
        (X"01",X"01",X"01",X"00",X"00",X"ba",X"ba",X"ba",X"ba",X"8c",X"8c",X"00",X"8c",X"00",X"01",X"01"),
        (X"01",X"01",X"00",X"9e",X"9e",X"2e",X"9e",X"ba",X"53",X"2e",X"00",X"8c",X"00",X"00",X"01",X"01"),
        (X"01",X"00",X"9e",X"9e",X"9e",X"9e",X"9e",X"9e",X"53",X"2e",X"00",X"00",X"8c",X"53",X"00",X"01"),
        (X"01",X"00",X"9e",X"2e",X"2e",X"9e",X"9e",X"9e",X"53",X"8c",X"8c",X"8c",X"8c",X"53",X"00",X"01"),
        (X"00",X"9e",X"9e",X"2e",X"2e",X"9e",X"9e",X"9e",X"9e",X"53",X"8c",X"8c",X"53",X"53",X"53",X"00"),
        (X"00",X"9e",X"9e",X"9e",X"9e",X"9e",X"9e",X"9e",X"9e",X"ba",X"53",X"53",X"53",X"53",X"53",X"00"),
        (X"00",X"9e",X"9e",X"9e",X"9e",X"9e",X"9e",X"9e",X"9e",X"ba",X"ba",X"ba",X"53",X"53",X"53",X"00"),
        (X"00",X"ba",X"9e",X"9e",X"9e",X"9e",X"9e",X"9e",X"ba",X"ba",X"ba",X"ba",X"53",X"53",X"53",X"00"),
        (X"00",X"ba",X"ba",X"9e",X"9e",X"9e",X"9e",X"ba",X"ba",X"ba",X"ba",X"53",X"53",X"53",X"53",X"00"),
        (X"00",X"53",X"ba",X"ba",X"ba",X"ba",X"ba",X"ba",X"ba",X"ba",X"ba",X"53",X"53",X"53",X"53",X"00"),
        (X"01",X"00",X"53",X"ba",X"ba",X"ba",X"ba",X"ba",X"ba",X"ba",X"53",X"53",X"53",X"53",X"00",X"01"),
        (X"01",X"00",X"53",X"53",X"ba",X"ba",X"ba",X"ba",X"53",X"53",X"53",X"53",X"53",X"53",X"00",X"01"),
        (X"01",X"01",X"00",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"00",X"01",X"01"),
        (X"01",X"01",X"01",X"00",X"00",X"53",X"53",X"53",X"53",X"53",X"53",X"00",X"00",X"01",X"01",X"01"),
        (X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01"));
end package;