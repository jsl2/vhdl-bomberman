library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

use work.graphics_pkg.all;
use work.touch_pkg.all;
use work.tileset_pkg.all;
use work.levels_pkg.all;
use work.maps_pkg.all;
use work.bombs_pkg.all;
use work.explosions_pkg.all;

package tile_state_pkg is  
    subtype tile_address is std_logic_vector(9 downto 0);
    
        type powerup_type is (bomb, blast, speed);
    type explosion_state_vector is record
        ACTIVE : boolean;
        FRAME : integer range 0 to 12; -- 4 bit
        DIR : direction;                -- 2 bit
        ORIG : boolean;
        EDGE : boolean;
        GOTO_NEXT_FRAME : boolean; -- toggle true false, i.e. slow animation
    end record; -- = 10 bit
    
    constant INITIAL_EXPLOSION_STATE : explosion_state_vector :=
        (ACTIVE => false,
         FRAME => 0,
         DIR => left,
         ORIG => false,
         EDGE => false,
         GOTO_NEXT_FRAME => false);
        
    
    type bomb_state_vector is record
        ACTIVE : boolean;
        FRAME : integer range 0 to 9; -- 4 bit
        COUNTER : integer range 0 to 23; -- 5 bit
    end record; -- = 10 bit
    
    constant INITIAL_BOMB_STATE : bomb_state_vector :=
        (ACTIVE => false,
         FRAME => 0,
         COUNTER => 0);
    
    type wall_state_vector is record
        ACTIVE : boolean;
        CRUMBLING : boolean;
        FRAME : integer range 0 to 7; --3 bit
        COUNTER : integer range 0 to 15; -- 4 bit
    end record; -- = 9 bit
    
    constant INITIAL_WALL_STATE : wall_state_vector :=
        (ACTIVE => false,
         CRUMBLING => false,
         FRAME => 0,
         COUNTER => 0);
    
    type powerup_state_vector is record
        ACTIVE : boolean;
        POWERUP_TYPE : powerup_type; -- 3 bit
    end record; -- 4 bit        
    
    constant INITIAL_POWERUP_STATE : powerup_state_vector :=
        (ACTIVE => false,
         POWERUP_TYPE => bomb);
    
    type tile_state_vector is record
        EXPLOSION : explosion_state_vector;
        BOMB : bomb_state_vector;
        WALL : wall_state_vector;
        POWERUP : powerup_state_vector;
    end record;
    
    constant INITIAL_TILE_STATE : tile_state_vector :=
        (EXPLOSION => INITIAL_EXPLOSION_STATE,
         BOMB => INITIAL_BOMB_STATE,
         WALL => INITIAL_WALL_STATE,
         POWERUP => INITIAL_POWERUP_STATE);
    
    subtype tile_state_slv is std_logic_vector(32 downto 0);
    type tile_state_ram is array (0 to 1023) of tile_state_slv;
    
    constant LEVEL0_STATE_RAM : tile_state_ram := 
    ('0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"60100000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"20100000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"20100000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"20100000",
    '0'&X"00100000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00100000",
    '0'&X"60100000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00100000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00100000",
    '0'&X"00100000",
    '0'&X"00100000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000",
    '0'&X"00000000");


    
    function pack_tile_state(in_state : in tile_state_vector) return tile_state_slv;
    function unpack_tile_state(in_state : in tile_state_slv) return tile_state_vector;      
end package;

package body tile_state_pkg is
        function pack_tile_state(in_state : in tile_state_vector) return tile_state_slv is
    variable ret : tile_state_slv:= (others => '0');
    variable current_bit : integer range 0 to 35 := 0;
begin
    current_bit := 0;
    if in_state.EXPLOSION.ACTIVE then
        ret(current_bit) := '1';
    else
        ret(current_bit) := '0';
    end if;        
    current_bit := current_bit + 1;
       
    ret(current_bit + 3 downto current_bit) := std_logic_vector(to_unsigned(in_state.EXPLOSION.FRAME,4));
    current_bit := current_bit + 4;
    
    case in_state.EXPLOSION.DIR is
        when left =>
            ret(current_bit+1 downto current_bit) := "00";
        when up =>
            ret(current_bit+1 downto current_bit) := "01";
        when right =>
            ret(current_bit+1 downto current_bit) := "10";
        when down =>
            ret(current_bit+1 downto current_bit) := "11";
    end case;
    current_bit := current_bit + 2;
    
    if in_state.EXPLOSION.ORIG then
        ret(current_bit) := '1';
    else
        ret(current_bit) := '0';
    end if;
    current_bit := current_bit + 1;                                                                  
    
    if in_state.EXPLOSION.EDGE then
        ret(current_bit) := '1';
    else
        ret(current_bit) := '0';
    end if;
    current_bit := current_bit + 1;
    
    if in_state.EXPLOSION.GOTO_NEXT_FRAME then
        ret(current_bit) := '1';
    else
        ret(current_bit) := '0';
    end if;
    current_bit := current_bit + 1;
    
    if in_state.BOMB.ACTIVE then
        ret(current_bit) := '1';
    else
        ret(current_bit) := '0';
    end if;
    current_bit := current_bit + 1;
    
    ret(current_bit + 3 downto current_bit) := std_logic_vector(to_unsigned(in_state.BOMB.FRAME,4));
    current_bit := current_bit + 4;
    
    ret(current_bit + 4 downto current_bit) := std_logic_vector(to_unsigned(in_state.BOMB.COUNTER,5));
    current_bit := current_bit + 5;
    
    if in_state.WALL.ACTIVE then
        ret(current_bit) := '1';
    else
        ret(current_bit) := '0';
    end if;
    current_bit := current_bit + 1;
    
    if in_state.WALL.CRUMBLING then
        ret(current_bit) := '1';
    else
        ret(current_bit) := '0';
    end if;
    current_bit := current_bit + 1;
    
    ret(current_bit + 2 downto current_bit) := std_logic_vector(to_unsigned(in_state.WALL.FRAME,3));
    current_bit := current_bit + 3;
    
    ret(current_bit + 3 downto current_bit) := std_logic_vector(to_unsigned(in_state.WALL.COUNTER,4));
    current_bit := current_bit + 4;
    
    if in_state.POWERUP.ACTIVE then
        ret(current_bit) := '1';
    else
        ret(current_bit) := '0';
    end if;        
    current_bit := current_bit + 1;
    
    case in_state.POWERUP.POWERUP_TYPE is
        when bomb =>
            ret(current_bit+2 downto current_bit) := "000";
        when blast =>
            ret(current_bit+2 downto current_bit) := "001";
        when speed =>
            ret(current_bit+2 downto current_bit) := "010";
        when others =>
            ret(current_bit+2 downto current_bit) := "111";
    end case;
    
    return ret;
end;

function unpack_tile_state(in_state : in tile_state_slv) return tile_state_vector is
    variable ret : tile_state_vector := INITIAL_TILE_STATE;
    variable current_bit : integer range 0 to 35 := 0;
begin
    current_bit := 0;
    
    ret.EXPLOSION.ACTIVE := in_state(current_bit) = '1';   
    current_bit := current_bit + 1;
    
    ret.EXPLOSION.FRAME := to_integer(unsigned(in_state(current_bit + 3 downto current_bit)));
    current_bit := current_bit + 4;
    
    case in_state(current_bit+1 downto current_bit) is
        when "00" =>
            ret.EXPLOSION.DIR := left;
        when "01" =>
            ret.EXPLOSION.DIR := up;
        when "10" =>
            ret.EXPLOSION.DIR := right;
        when "11" =>
            ret.EXPLOSION.DIR := down;
    end case;
    current_bit := current_bit + 2;
    
    ret.EXPLOSION.ORIG := in_state(current_bit) = '1';   
    current_bit := current_bit + 1;                                                               

    ret.EXPLOSION.EDGE := in_state(current_bit) = '1';   
    current_bit := current_bit + 1;        
    
    ret.EXPLOSION.GOTO_NEXT_FRAME := in_state(current_bit) = '1';   
    current_bit := current_bit + 1;        
    
    ret.BOMB.ACTIVE := in_state(current_bit) = '1';   
    current_bit := current_bit + 1;        

    ret.BOMB.FRAME := to_integer(unsigned(in_state(current_bit + 3 downto current_bit)));
    current_bit := current_bit + 4;

    ret.BOMB.COUNTER := to_integer(unsigned(in_state(current_bit + 4 downto current_bit)));
    current_bit := current_bit + 5;       

    ret.WALL.ACTIVE := in_state(current_bit) = '1';   
    current_bit := current_bit + 1;        

    ret.WALL.CRUMBLING := in_state(current_bit) = '1';   
    current_bit := current_bit + 1;
           
    ret.WALL.FRAME := to_integer(unsigned(in_state(current_bit + 2 downto current_bit)));
    current_bit := current_bit + 3;       
    
    ret.WALL.COUNTER := to_integer(unsigned(in_state(current_bit + 3 downto current_bit)));
    current_bit := current_bit + 4;                

    ret.POWERUP.ACTIVE  := in_state(current_bit) = '1';   
    current_bit := current_bit + 1;        
    
    case in_state(current_bit+2 downto current_bit) is
        when "000" =>
            ret.POWERUP.POWERUP_TYPE := bomb;
        when "001" =>
            ret.POWERUP.POWERUP_TYPE := blast;
        when "010" =>
            ret.POWERUP.POWERUP_TYPE := speed;
        when others =>
            ret.POWERUP.POWERUP_TYPE := bomb;
            ret.POWERUP.ACTIVE := false;
    end case;
    
    return ret;
end;
end; 